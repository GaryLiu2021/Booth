
module booth_multiplier (multiplicand, multiplier, result);
 input [31:0] multiplicand;
 input [31:0] multiplier;
 output [63:0] result;
  wire VCC_NET;
  wire GND_NET;
  wire id02400;
  wire id02401;
  wire id02402;
  wire id02403;
  wire id02404;
  wire id02405;
  wire id02406;
  wire id02407;
  wire id02408;
  wire id02409;
  wire id02410;
  wire id02411;
  wire id02412;
  wire id02413;
  wire id02414;
  wire id02415;
  wire id02416;
  wire id02417;
  wire id02418;
  wire id02419;
  wire id02420;
  wire id02421;
  wire id02422;
  wire id02423;
  wire id02424;
  wire id02425;
  wire id02426;
  wire id02427;
  wire id02428;
  wire id02429;
  wire id02430;
  wire id02431;
  wire id02432;
  wire id02433;
  wire id02434;
  wire id02435;
  wire id02436;
  wire id02437;
  wire id02438;
  wire id02439;
  wire id02440;
  wire id02441;
  wire \u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ;
  wire id02444;
  wire id02445;
  wire id02446;
  wire id02447;
  wire \u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[40].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 ;
  wire id02452;
  wire id02453;
  wire id02454;
  wire id02455;
  wire id02456;
  wire id02457;
  wire id02458;
  wire id02459;
  wire id02460;
  wire id02461;
  wire id02462;
  wire id02463;
  wire id02464;
  wire id02465;
  wire id02466;
  wire id02467;
  wire id02468;
  wire id02469;
  wire id02470;
  wire id02471;
  wire id02472;
  wire id02473;
  wire id02474;
  wire id02475;
  wire id02476;
  wire id02477;
  wire id02478;
  wire id02479;
  wire id02480;
  wire id02481;
  wire id02482;
  wire id02483;
  wire id02484;
  wire id02485;
  wire id02486;
  wire id02487;
  wire id02488;
  wire id02489;
  wire id02490;
  wire id02491;
  wire id02492;
  wire id02493;
  wire id02494;
  wire id02495;
  wire id02496;
  wire id02497;
  wire id02498;
  wire id02499;
  wire id02500;
  wire id02501;
  wire id02502;
  wire id02503;
  wire id02504;
  wire id02505;
  wire id02506;
  wire id02507;
  wire id02508;
  wire id02509;
  wire id02510;
  wire id02511;
  wire id02512;
  wire id02513;
  wire id02514;
  wire id02515;
  wire id02516;
  wire id02517;
  wire id02518;
  wire id02519;
  wire id02520;
  wire \u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[40].u_compressor42_cell.x3 ;
  wire id02523;
  wire id02524;
  wire id02525;
  wire id02526;
  wire id02527;
  wire id02528;
  wire id02529;
  wire id02530;
  wire id02531;
  wire id02532;
  wire id02533;
  wire id02534;
  wire id02535;
  wire id02536;
  wire id02537;
  wire id02538;
  wire id02539;
  wire id02540;
  wire id02541;
  wire id02542;
  wire id02543;
  wire id02544;
  wire id02545;
  wire id02546;
  wire id02547;
  wire id02548;
  wire id02549;
  wire id02550;
  wire id02551;
  wire id02552;
  wire id02553;
  wire id02554;
  wire id02555;
  wire id02556;
  wire id02557;
  wire id02558;
  wire id02559;
  wire id02560;
  wire id02561;
  wire id02562;
  wire id02563;
  wire id02564;
  wire id02565;
  wire id02566;
  wire id02567;
  wire id02568;
  wire id02569;
  wire id02570;
  wire id02571;
  wire id02572;
  wire id02573;
  wire id02574;
  wire id02575;
  wire id02576;
  wire id02577;
  wire id02578;
  wire id02579;
  wire id02580;
  wire id02581;
  wire id02582;
  wire id02583;
  wire id02584;
  wire id02585;
  wire id02586;
  wire id02587;
  wire id02588;
  wire id02589;
  wire id02590;
  wire id02591;
  wire id02592;
  wire id02593;
  wire id02594;
  wire id02595;
  wire id02596;
  wire id02597;
  wire \u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[39].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[2].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 ;
  wire id02683;
  wire id02684;
  wire id02685;
  wire id02686;
  wire id02687;
  wire id02688;
  wire id02689;
  wire id02690;
  wire id02691;
  wire id02692;
  wire id02693;
  wire id02694;
  wire id02695;
  wire id02696;
  wire id02697;
  wire id02698;
  wire id02699;
  wire \u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[38].u_compressor42_cell.x3 ;
  wire id02703;
  wire \u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 ;
  wire id02705;
  wire id02706;
  wire id02707;
  wire id02708;
  wire id02709;
  wire id02710;
  wire \u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x0 ;
  wire id02758;
  wire id02759;
  wire id02760;
  wire id02761;
  wire id02762;
  wire id02763;
  wire id02764;
  wire id02765;
  wire id02766;
  wire id02767;
  wire id02768;
  wire id02769;
  wire id02770;
  wire id02771;
  wire id02772;
  wire id02773;
  wire id02774;
  wire id02775;
  wire id02776;
  wire id02777;
  wire id02778;
  wire id02779;
  wire id02780;
  wire id02781;
  wire id02782;
  wire id02783;
  wire id02784;
  wire id02785;
  wire id02786;
  wire id02787;
  wire id02788;
  wire id02789;
  wire id02790;
  wire id02791;
  wire id02792;
  wire id02793;
  wire id02794;
  wire id02795;
  wire id02796;
  wire id02797;
  wire id02798;
  wire id02799;
  wire id02800;
  wire id02801;
  wire id02802;
  wire id02803;
  wire id02804;
  wire id02805;
  wire id02806;
  wire id02807;
  wire id02808;
  wire id02809;
  wire id02810;
  wire id02811;
  wire id02812;
  wire id02813;
  wire id02814;
  wire id02815;
  wire id02816;
  wire id02817;
  wire id02818;
  wire id02819;
  wire id02820;
  wire id02821;
  wire id02822;
  wire id02823;
  wire id02824;
  wire id02825;
  wire id02826;
  wire id02827;
  wire id02828;
  wire id02829;
  wire id02830;
  wire id02831;
  wire \u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[2].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x2 ;
  wire id02978;
  wire id02979;
  wire \u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[2].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x3 ;
  wire id03085;
  wire id03086;
  wire \u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x0 ;
  wire \DECODE_GEN[3].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[7].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[6].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[5].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[4].u_booth_enc.partial_reverse ;
  wire id03154;
  wire id03155;
  wire id03156;
  wire id03157;
  wire id03158;
  wire id03159;
  wire id03160;
  wire id03161;
  wire id03162;
  wire id03163;
  wire id03164;
  wire id03165;
  wire id03166;
  wire id03167;
  wire id03168;
  wire id03169;
  wire id03170;
  wire id03171;
  wire id03172;
  wire id03173;
  wire id03174;
  wire id03175;
  wire id03176;
  wire id03177;
  wire id03178;
  wire id03179;
  wire id03180;
  wire id03181;
  wire id03182;
  wire id03183;
  wire id03184;
  wire id03185;
  wire id03186;
  wire id03187;
  wire id03188;
  wire id03189;
  wire id03190;
  wire id03191;
  wire id03192;
  wire id03193;
  wire id03194;
  wire id03195;
  wire id03196;
  wire id03197;
  wire id03198;
  wire id03199;
  wire id03200;
  wire id03201;
  wire id03202;
  wire id03203;
  wire id03204;
  wire id03205;
  wire id03206;
  wire id03207;
  wire id03208;
  wire id03209;
  wire id03210;
  wire id03211;
  wire id03212;
  wire id03213;
  wire id03214;
  wire id03215;
  wire id03216;
  wire id03217;
  wire id03218;
  wire id03219;
  wire id03220;
  wire id03221;
  wire id03222;
  wire id03223;
  wire id03224;
  wire id03225;
  wire id03226;
  wire id03227;
  wire id03228;
  wire id03229;
  wire id03230;
  wire id03231;
  wire id03232;
  wire id03233;
  wire id03234;
  wire id03235;
  wire id03236;
  wire id03237;
  wire id03238;
  wire id03239;
  wire id03240;
  wire id03241;
  wire id03242;
  wire id03243;
  wire id03244;
  wire id03245;
  wire id03246;
  wire id03247;
  wire id03248;
  wire id03249;
  wire id03250;
  wire id03251;
  wire id03252;
  wire id03253;
  wire id03254;
  wire id03255;
  wire id03256;
  wire id03257;
  wire id03258;
  wire id03259;
  wire id03260;
  wire id03261;
  wire id03262;
  wire id03263;
  wire id03264;
  wire id03265;
  wire id03266;
  wire id03267;
  wire id03268;
  wire id03269;
  wire id03270;
  wire id03271;
  wire id03272;
  wire id03273;
  wire id03274;
  wire id03275;
  wire id03276;
  wire id03277;
  wire id03278;
  wire id03279;
  wire \net_Buf-pad-multiplicand[16] ;
  wire \net_Buf-pad-multiplicand[17] ;
  wire \net_Buf-pad-multiplicand[18] ;
  wire \net_Buf-pad-multiplicand[19] ;
  wire \net_Buf-pad-multiplicand[20] ;
  wire \net_Buf-pad-multiplicand[21] ;
  wire \net_Buf-pad-multiplicand[22] ;
  wire \net_Buf-pad-multiplicand[23] ;
  wire \net_Buf-pad-multiplicand[24] ;
  wire \net_Buf-pad-multiplicand[25] ;
  wire \net_Buf-pad-multiplicand[26] ;
  wire \net_Buf-pad-multiplicand[27] ;
  wire \net_Buf-pad-multiplicand[28] ;
  wire \net_Buf-pad-multiplicand[29] ;
  wire \net_Buf-pad-multiplicand[30] ;
  wire \net_Buf-pad-multiplicand[31] ;
  wire \net_Buf-pad-multiplicand[0] ;
  wire \net_Buf-pad-multiplicand[1] ;
  wire \net_Buf-pad-multiplicand[2] ;
  wire \net_Buf-pad-multiplicand[3] ;
  wire \net_Buf-pad-multiplicand[4] ;
  wire \net_Buf-pad-multiplicand[5] ;
  wire \net_Buf-pad-multiplicand[6] ;
  wire \net_Buf-pad-multiplicand[7] ;
  wire \net_Buf-pad-multiplicand[8] ;
  wire \net_Buf-pad-multiplicand[9] ;
  wire \net_Buf-pad-multiplicand[10] ;
  wire \net_Buf-pad-multiplicand[11] ;
  wire \net_Buf-pad-multiplicand[12] ;
  wire \net_Buf-pad-multiplicand[13] ;
  wire \net_Buf-pad-multiplicand[14] ;
  wire \net_Buf-pad-multiplicand[15] ;
  wire id03312;
  wire \net_Buf-pad-result[18] ;
  wire \net_Buf-pad-result[19] ;
  wire \net_Buf-pad-result[16] ;
  wire \net_Buf-pad-result[17] ;
  wire \net_Buf-pad-result[22] ;
  wire \net_Buf-pad-result[23] ;
  wire \net_Buf-pad-result[20] ;
  wire \net_Buf-pad-result[21] ;
  wire \net_Buf-pad-result[26] ;
  wire \net_Buf-pad-result[27] ;
  wire \net_Buf-pad-result[24] ;
  wire \net_Buf-pad-result[25] ;
  wire \net_Buf-pad-result[30] ;
  wire \net_Buf-pad-result[31] ;
  wire \net_Buf-pad-result[28] ;
  wire \net_Buf-pad-result[29] ;
  wire \net_Buf-pad-result[6] ;
  wire \net_Buf-pad-result[7] ;
  wire \net_Buf-pad-result[4] ;
  wire \net_Buf-pad-result[5] ;
  wire \net_Buf-pad-result[10] ;
  wire \net_Buf-pad-result[11] ;
  wire \net_Buf-pad-result[8] ;
  wire \net_Buf-pad-result[9] ;
  wire \net_Buf-pad-result[14] ;
  wire \net_Buf-pad-result[15] ;
  wire \net_Buf-pad-result[12] ;
  wire \net_Buf-pad-result[13] ;
  wire \net_Buf-pad-multiplier[19] ;
  wire \net_Buf-pad-result[50] ;
  wire \net_Buf-pad-multiplier[18] ;
  wire \net_Buf-pad-result[51] ;
  wire \net_Buf-pad-multiplier[17] ;
  wire \net_Buf-pad-result[48] ;
  wire \net_Buf-pad-multiplier[16] ;
  wire \net_Buf-pad-result[49] ;
  wire \net_Buf-pad-multiplier[23] ;
  wire \net_Buf-pad-result[54] ;
  wire \net_Buf-pad-multiplier[22] ;
  wire \net_Buf-pad-result[55] ;
  wire \net_Buf-pad-multiplier[21] ;
  wire \net_Buf-pad-result[52] ;
  wire \net_Buf-pad-multiplier[20] ;
  wire \net_Buf-pad-result[53] ;
  wire \net_Buf-pad-multiplier[27] ;
  wire \net_Buf-pad-result[58] ;
  wire \net_Buf-pad-multiplier[26] ;
  wire \net_Buf-pad-result[59] ;
  wire \net_Buf-pad-multiplier[25] ;
  wire \net_Buf-pad-result[56] ;
  wire \net_Buf-pad-multiplier[24] ;
  wire \net_Buf-pad-result[57] ;
  wire \net_Buf-pad-multiplier[31] ;
  wire \net_Buf-pad-result[62] ;
  wire \net_Buf-pad-multiplier[30] ;
  wire \net_Buf-pad-result[63] ;
  wire \net_Buf-pad-multiplier[29] ;
  wire \net_Buf-pad-result[60] ;
  wire \net_Buf-pad-multiplier[28] ;
  wire \net_Buf-pad-result[61] ;
  wire \net_Buf-pad-multiplier[3] ;
  wire \net_Buf-pad-result[34] ;
  wire \net_Buf-pad-multiplier[2] ;
  wire \net_Buf-pad-result[35] ;
  wire \net_Buf-pad-multiplier[1] ;
  wire \net_Buf-pad-result[32] ;
  wire \net_Buf-pad-multiplier[0] ;
  wire \net_Buf-pad-result[33] ;
  wire \net_Buf-pad-multiplier[7] ;
  wire \net_Buf-pad-result[38] ;
  wire \net_Buf-pad-multiplier[6] ;
  wire \net_Buf-pad-result[39] ;
  wire \net_Buf-pad-multiplier[5] ;
  wire \net_Buf-pad-result[36] ;
  wire \net_Buf-pad-multiplier[4] ;
  wire \net_Buf-pad-result[37] ;
  wire \net_Buf-pad-multiplier[11] ;
  wire \net_Buf-pad-result[42] ;
  wire \net_Buf-pad-multiplier[10] ;
  wire \net_Buf-pad-result[43] ;
  wire \net_Buf-pad-multiplier[9] ;
  wire \net_Buf-pad-result[40] ;
  wire \net_Buf-pad-multiplier[8] ;
  wire \net_Buf-pad-result[41] ;
  wire \net_Buf-pad-multiplier[15] ;
  wire \net_Buf-pad-result[46] ;
  wire \net_Buf-pad-multiplier[14] ;
  wire \net_Buf-pad-result[47] ;
  wire \net_Buf-pad-multiplier[13] ;
  wire \net_Buf-pad-result[44] ;
  wire \net_Buf-pad-multiplier[12] ;
  wire \net_Buf-pad-result[45] ;
  wire id03405;
  wire id03406;
  wire id03407;
  wire id03408;
  wire id03409;
  wire id03410;
  wire id03411;
  wire id03412;
  wire id03413;
  wire \DECODE_GEN[2].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[1].u_booth_enc.partial_reverse ;
  wire id03416;
  wire id03417;
  wire id03418;
  wire id03419;
  wire id03420;
  wire id03421;
  wire id03422;
  wire id03423;
  wire id03424;
  wire id03425;
  wire id03426;
  wire id03427;
  wire id03428;
  wire id03429;
  wire id03430;
  wire id03431;
  wire id03432;
  wire id03433;
  wire id03434;
  wire id03435;
  wire id03436;
  wire id03437;
  wire id03438;
  wire id03439;
  wire id03440;
  wire id03441;
  wire id03442;
  wire id03443;
  wire id03444;
  wire id03445;
  wire id03446;
  wire id03447;
  wire id03448;
  wire id03449;
  wire id03450;
  wire id03451;
  wire id03452;
  wire id03453;
  wire id03454;
  wire id03455;
  wire id03456;
  wire id03457;
  wire id03458;
  wire id03459;
  wire id03460;
  wire id03461;
  wire id03462;
  wire id03463;
  wire id03464;
  wire id03465;
  wire id03466;
  wire id03467;
  wire id03468;
  wire id03469;
  wire id03470;
  wire id03471;
  wire id03472;
  wire id03473;
  wire id03474;
  wire id03475;
  wire id03476;
  wire id03477;
  wire id03478;
  wire id03479;
  wire id03480;
  wire id03481;
  wire id03482;
  wire id03483;
  wire id03484;
  wire id03485;
  wire id03486;
  wire id03487;
  wire id03488;
  wire id03489;
  wire id03490;
  wire id03491;
  wire id03492;
  wire id03493;
  wire id03494;
  wire id03495;
  wire id03496;
  wire id03497;
  wire id03498;
  wire id03499;
  wire id03500;
  wire id03501;
  wire id03502;
  wire id03503;
  wire id03504;
  wire id03505;
  wire id03506;
  wire id03507;
  wire id03508;
  wire id03509;
  wire id03510;
  wire id03511;
  wire id03512;
  wire id03513;
  wire id03514;
  wire id03515;
  wire id03516;
  wire id03517;
  wire id03518;
  wire id03519;
  wire id03520;
  wire id03521;
  wire id03522;
  wire id03523;
  wire id03524;
  wire id03525;
  wire id03526;
  wire id03527;
  wire id03528;
  wire id03529;
  wire id03530;
  wire id03531;
  wire id03532;
  wire id03533;
  wire id03534;
  wire id03535;
  wire id03536;
  wire id03537;
  wire id03538;
  wire id03539;
  wire id03540;
  wire id03541;
  wire id03542;
  wire id03543;
  wire id03544;
  wire id03545;
  wire id03546;
  wire id03547;
  wire id03548;
  wire id03549;
  wire id03550;
  wire id03551;
  wire id03552;
  wire id03553;
  wire id03554;
  wire id03555;
  wire id03556;
  wire id03557;
  wire id03558;
  wire id03559;
  wire id03560;
  wire id03561;
  wire id03562;
  wire id03563;
  wire id03564;
  wire id03565;
  wire id03566;
  wire id03567;
  wire id03568;
  wire id03569;
  wire id03570;
  wire id03571;
  wire id03572;
  wire id03573;
  wire id03574;
  wire id03575;
  wire id03576;
  wire id03577;
  wire id03578;
  wire id03579;
  wire id03580;
  wire id03581;
  wire id03582;
  wire id03583;
  wire id03584;
  wire id03585;
  wire id03586;
  wire id03587;
  wire id03588;
  wire id03589;
  wire id03590;
  wire id03591;
  wire id03592;
  wire id03593;
  wire id03594;
  wire id03595;
  wire id03596;
  wire id03597;
  wire id03598;
  wire id03599;
  wire id03600;
  wire id03601;
  wire id03602;
  wire id03603;
  wire id03604;
  wire id03605;
  wire id03606;
  wire id03607;
  wire id03608;
  wire \u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x1 ;
  wire id03621;
  wire id03622;
  wire id03623;
  wire id03624;
  wire \u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x0 ;
  wire id03632;
  wire id03633;
  wire id03634;
  wire id03635;
  wire id03636;
  wire id03637;
  wire id03638;
  wire id03639;
  wire \u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 ;
  wire id03641;
  wire id03642;
  wire \u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x0 ;
  wire id03645;
  wire \u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x1 ;
  wire id03647;
  wire \u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x0 ;
  wire id03649;
  wire id03650;
  wire id03651;
  wire id03652;
  wire id03653;
  wire \u_compressor42_l0_0.CELLS[0].u_compressor42_cell.x0 ;
  wire id03655;
  wire id03656;
  wire id03657;
  wire id03658;
  wire \u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x2 ;
  wire \u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x1 ;
  wire \u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x0 ;
  wire \u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x3 ;
  wire \u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x2 ;
  wire \DECODE_GEN[11].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[10].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[9].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[8].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[14].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[13].u_booth_enc.partial_reverse ;
  wire \DECODE_GEN[12].u_booth_enc.partial_reverse ;
  wire id03713;
  wire id03714;
  wire id03715;
  wire id03716;
  wire id03717;
  wire id03718;
  wire id03719;
  wire id03720;
  wire id03721;
  wire id03722;
  wire id03723;
  wire id03724;
  wire id03725;
  wire id03726;
  wire id03727;
  wire id03728;
  wire id03729;
  wire id03730;
  wire id03731;
  wire id03732;
  wire id03733;
  wire id03734;
  wire id03735;
  wire id03736;
  wire id03737;
  wire id03738;
  wire id03739;
  wire id03740;
  wire id03741;
  wire id03742;
  wire id03743;
  wire id03744;
  wire id03745;
  wire id03746;
  wire id03747;
  wire id03748;
  wire id03749;
  wire id03750;
  wire id03751;
  wire id03752;
  wire id03753;
  wire id03754;
  wire id03755;
  wire id03756;
  wire id03757;
  wire id03758;
  wire id03759;
  wire id03760;
  wire id03761;
  wire id03762;
  wire id03763;
  wire id03764;
  wire id03765;
  wire id03766;
  wire id03767;
  wire id03768;
  wire id03769;
  wire id03770;
  wire id03771;
  wire id03772;
  wire id03773;
  wire id03774;
  wire id03775;
  wire id03776;
  wire id03777;
  wire id03778;
  wire id03779;
  wire id03780;
  wire id03781;
  wire id03782;
  wire id03783;
  wire id03784;
  wire id03785;
  wire id03786;
  wire id03787;
  wire id03788;
  wire id03789;
  wire id03790;
  wire id03791;
  wire id03792;
  wire id03793;
  wire id03794;
  wire id03795;
  wire id03796;
  wire id03797;
  wire id03798;
  wire id03799;
  wire id03800;
  wire id03801;
  wire id03802;
  wire id03803;
  wire id03804;
  wire id03805;
  wire id03806;
  wire id03807;
  wire id03808;
  wire id03809;
  wire id03810;
  wire id03811;
  wire id03812;
  wire id03813;
  wire id03814;
  wire id03815;
  wire id03816;
  wire id03817;
  wire id03818;
  wire id03819;
  wire id03820;
  wire id03821;
  wire id03822;
  wire id03823;
  wire id03824;
  wire id03825;
  wire id03826;
  wire id03827;
  wire id03828;
  wire id03829;
  wire id03830;
  wire id03831;
  wire id03832;
  wire id03833;
  wire id03834;
  wire id03835;
  wire id03836;
  wire id03837;
  wire id03838;
  wire id03839;
  wire id03840;
  wire id03841;
  wire id03842;
  wire id03843;
  wire id03844;
  wire id03845;
  wire id03846;
  wire id03847;
  wire id03848;
  wire id03849;
  wire id03850;
  wire id03851;
  wire id03852;
  wire id03853;
  wire id03854;
  wire id03855;
  wire id03856;
  wire id03857;
  wire id03858;
  wire id03859;
  wire id03860;
  wire id03861;
  wire id03862;
  wire id03863;
  wire id03864;
  wire id03865;
  wire id03866;
  wire id03867;
  wire id03868;
  wire id03869;
  wire id03870;
  wire id03871;
  wire id03872;
  wire id03873;
  wire id03874;
  wire id03875;
  wire id03876;
  wire id03877;
  wire id03878;
  wire id03879;
  wire id03880;
  wire id03881;
  wire id03882;
  wire id03883;
  wire id03884;
  wire id03885;
  wire id03886;
  wire id03887;
  wire id03888;
  wire id03889;
  wire id03890;
  wire id03891;
  wire id03892;
  wire id03893;
  wire id03894;
  wire id03895;
  wire id03896;
  wire id03897;
  wire id03898;
  wire id03899;
  wire id03900;
  wire id03901;
  wire id03902;
  wire id03903;
  wire id03904;
  wire id03905;
  wire id03906;
  wire id03907;
  wire id03908;
  wire id03909;
  wire id03910;
  wire id03911;
  wire id03912;
  wire id03913;
  wire id03914;
  wire id03915;
  wire id03916;
  wire id03917;
  wire id03918;
  wire id03919;
  wire id03920;
  wire id03921;
  wire id03922;
  wire id03923;
  wire id03924;
  wire id03925;
  wire id03926;
  wire id03927;
  wire id03928;
  wire id03929;
  wire id03930;
  wire id03931;
  wire id03932;
  wire id03933;
  wire id03934;
  wire id03935;
  wire id03936;
  wire id03937;
  wire id03938;
  wire id03939;
  wire id03940;
  wire id03941;
  wire id03942;
  wire id03943;
  wire id03944;
  wire id03945;
  wire id03946;
  wire id03947;
  wire id03948;
  wire id03949;
  wire id03950;
  wire id03951;
  wire id03952;
  wire id03953;
  wire id03954;
  wire id03955;
  wire id03956;
  wire id03957;
  wire id03958;
  wire id03959;
  wire id03960;
  wire id03961;
  wire id03962;
  wire id03963;
  wire id03964;
  wire id03965;
  wire id03966;
  wire id03967;
  wire id03968;
  wire id03969;
  wire id03970;
  wire id03971;
  wire id03972;
  wire id03973;
  wire id03974;
  wire id03975;
  wire id03976;
  wire id03977;
  wire id03978;
  wire id03979;
  wire id03980;
  wire id03981;
  wire id03982;
  wire id03983;
  wire id03984;
  wire id03985;
  wire id03986;
  wire id03987;
  wire id03988;
  wire id03989;
  wire id03990;
  wire id03991;
  wire id03992;
  wire id03993;
  wire id03994;
  wire id03995;
  wire id03996;
  wire id03997;
  wire id03998;
  wire id03999;
  wire id04000;
  wire id04001;
  wire id04002;
  wire id04003;
  wire id04004;
  wire id04005;
  wire id04006;
  wire id04007;
  wire id04008;
  wire id04009;
  wire id04010;
  wire id04011;
  wire id04012;
  wire id04013;
  wire id04014;
  wire id04015;
  wire id04016;
  wire id04017;
  wire id04018;
  wire id04019;
  wire id04020;
  wire id04021;
  wire id04022;
  wire id04023;
  wire id04024;
  wire id04025;
  wire id04026;
  wire id04027;
  wire id04028;
  wire id04029;
  wire id04030;
  wire id04031;
  wire id04032;
  wire id04033;
  wire id04034;
  wire id04035;
  wire id04036;
  wire id04037;
  wire id04038;
  wire id04039;
  wire id04040;
  wire id04041;
  wire id04042;
  wire id04043;
  wire id04044;
  wire id04045;
  wire id04046;
  wire id04047;
  wire id04048;
  wire id04049;
  wire id04050;
  wire id04051;
  wire id04052;
  wire id04053;
  wire id04054;
  wire id04055;
  wire id04056;
  wire id04057;
  wire id04058;
  wire id04059;
  wire id04060;
  wire id04061;
  wire id04062;
  wire id04063;
  wire id04064;
  wire id04065;
  wire id04066;
  wire id04067;
  wire id04068;
  wire id04069;
  wire id04070;
  wire id04071;
  wire id04072;
  wire id04073;
  wire id04074;
  wire id04075;
  wire id04076;
  wire id04077;
  wire id04078;
  wire id04079;
  wire id04080;
  wire id04081;
  wire id04082;
  wire id04083;
  wire id04084;
  wire id04085;
  wire id04086;
  wire id04087;
  wire id04088;
  wire id04089;
  wire id04090;
  wire id04091;
  wire id04092;
  wire id04093;
  wire id04094;
  wire id04095;
  wire id04096;
  wire id04097;
  wire id04098;
  wire id04099;
  wire id04100;
  wire id04101;
  wire id04102;
  wire id04103;
  wire id04104;
  wire id04105;
  wire id04106;
  wire id04107;
  wire id04108;
  wire id04109;
  wire id04110;
  wire id04111;
  wire id04112;
  wire id04113;
  wire id04114;
  wire id04115;
  wire id04116;
  wire id04117;
  wire id04118;
  wire id04119;
  wire id04120;
  wire id04121;
  wire id04122;
  wire id04123;
  wire id04124;
  wire id04125;
  wire id04126;
  wire id04127;
  wire id04128;
  wire id04129;
  wire id04130;
  wire id04131;
  wire id04132;
  wire id04133;
  wire id04134;
  wire id04135;
  wire id04136;
  wire id04137;
  wire id04138;
  wire id04139;
  wire id04140;
  wire id04141;
  wire id04142;
  wire id04143;
  wire id04144;
  wire id04145;
  wire id04146;
  wire id04147;
  wire id04148;
  wire id04149;
  wire id04150;
  wire id04151;
  wire id04152;
  wire id04153;
  wire id04154;
  wire id04155;
  wire id04156;
  wire id04157;
  wire id04158;
  wire id04159;
  wire id04160;
  wire id04161;
  wire id04162;
  wire id04163;
  wire id04164;
  wire id04165;
  wire id04166;
  wire id04167;
  wire id04168;
  wire id04169;
  wire id04170;
  wire id04171;
  wire id04172;
  wire id04173;
  wire id04174;
  wire id04175;
  wire id04176;
  wire id04177;
  wire id04178;
  wire id04179;
  wire id04180;
  wire id04181;
  wire id04182;
  wire id04183;
  wire id04184;
  wire id04185;
  wire id04186;
  wire id04187;
  wire id04188;
  wire id04189;
  wire id04190;
  wire id04191;
  wire id04192;
  wire id04193;
  wire id04194;
  wire id04195;
  wire id04196;
  wire id04197;
  wire id04198;
  wire id04199;
  wire id04200;
  wire id04201;
  wire id04202;
  wire id04203;
  wire id04204;
  wire id04205;
  wire id04206;
  wire id04207;
  wire id04208;
  wire id04209;
  wire id04210;
  wire id04211;
  wire id04212;
  wire id04213;
  wire id04214;
  wire id04215;
  wire id04216;
  wire id04217;
  wire id04218;
  wire id04219;
  wire id04220;
  wire id04221;
  wire id04222;
  wire id04223;
  wire id04224;
  wire id04225;
  wire id04226;
  wire id04227;
  wire id04228;
  wire id04229;
  wire id04230;
  wire id04231;
  wire id04232;
  wire id04233;
  wire id04234;
  wire id04235;
  wire id04236;
  wire id04237;
  wire id04238;
  wire id04239;
  wire id04240;
  wire id04241;
  wire id04242;
  wire id04243;
  wire id04244;
  wire id04245;
  wire id04246;
  wire id04247;
  wire id04248;
  wire id04249;
  wire id04250;
  wire id04251;
  wire id04252;
  wire id04253;
  wire id04254;
  wire id04255;
  wire id04256;
  wire id04257;
  wire id04258;
  wire id04259;
  wire id04260;
  wire id04261;
  wire id04262;
  wire id04263;
  wire id04264;
  wire id04265;
  wire id04266;
  wire id04267;
  wire id04268;
  wire id04269;
  wire id04270;
  wire id04271;
  wire id04272;
  wire id04273;
  wire id04274;
  wire id04275;
  wire id04276;
  wire id04277;
  wire id04278;
  wire id04279;
  wire id04280;
  wire id04281;
  wire id04282;
  wire id04283;
  wire id04284;
  wire id04285;
  wire id04286;
  wire id04287;
  wire id04288;
  wire id04289;
  wire id04290;
  wire id04291;
  wire id04292;
  wire id04293;
  wire id04294;
  wire id04295;
  wire id04296;
  wire id04297;
  wire id04298;
  wire id04299;
  wire id04300;
  wire id04301;
  wire id04302;
  wire id04303;
  wire id04304;
  wire id04305;
  wire id04306;
  wire id04307;
  wire id04308;
  wire id04309;
  wire id04310;
  wire id04311;
  wire id04312;
  wire id04313;
  wire id04314;
  wire id04315;
  wire id04316;
  wire id04317;
  wire id04318;
  wire id04319;
  wire id04320;
  wire id04321;
  wire id04322;
  wire id04323;
  wire id04324;
  wire id04325;
  wire id04326;
  wire id04327;
  wire id04328;
  wire id04329;
  wire id04330;
  wire id04331;
  wire id04332;
  wire id04333;
  wire id04334;
  wire id04335;
  wire id04336;
  wire id04337;
  wire id04338;
  wire id04339;
  wire id04340;
  wire id04341;
  wire id04342;
  wire id04343;
  wire id04344;
  wire id04345;
  wire id04346;
  wire id04347;
  wire id04348;
  wire id04349;
  wire id04350;
  wire id04351;
  wire id04352;
  wire id04353;
  wire id04354;
  wire id04355;
  wire id04356;
  wire id04357;
  wire id04358;
  wire id04359;
  wire id04360;
  wire id04361;
  wire id04362;
  wire id04363;
  wire id04364;
  wire id04365;
  wire id04366;
  wire id04367;
  wire id04368;
  wire id04369;
  wire id04370;
  wire id04371;
  wire id04372;
  wire id04373;
  wire id04374;
  wire id04375;
  wire id04376;
  wire id04377;
  wire id04378;
  wire id04379;
  wire id04380;
  wire id04381;
  wire id04382;
  wire id04383;
  wire id04384;
  wire id04385;
  wire id04386;
  wire id04387;
  wire id04388;
  wire id04389;
  wire id04390;
  wire id04391;
  wire id04392;
  wire id04393;
  wire id04394;
  wire id04395;
  wire id04396;
  wire id04397;
  wire id04398;
  wire id04399;
  wire id04400;
  wire id04401;
  wire id04402;
  wire id04403;
  wire id04404;
  wire id04405;
  wire id04406;
  wire id04407;
  wire id04408;
  wire id04409;
  wire id04410;
  wire id04411;
  wire id04412;
  wire id04413;
  wire id04414;
  wire id04415;
  wire id04416;
  wire id04417;
  wire id04418;
  wire id04419;
  wire id04420;
  wire id04421;
  wire id04422;
  wire id04423;
  wire id04424;
  wire id04425;
  wire id04426;
  wire id04427;
  wire id04428;
  wire id04429;
  wire id04430;
  wire id04431;
  wire id04432;
  wire id04433;
  wire id04434;
  wire id04435;
  wire id04436;
  wire id04437;
  wire id04438;
  wire id04439;
  wire id04440;
  wire id04441;
  wire id04442;
  wire id04443;
  wire id04444;
  wire id04445;
  wire id04446;
  wire id04447;
  wire id04448;
  wire id04449;
  wire id04450;
  wire id04451;
  wire id04452;
  wire id04453;
  wire id04454;
  wire id04455;
  wire id04456;
  wire id04457;
  wire id04458;
  wire id04459;
  wire id04460;
  wire id04461;
  wire id04462;
  wire id04463;
  wire id04464;
  wire id04465;
  wire id04466;
  wire id04467;
  wire id04468;
  wire id04469;
  wire id04470;
  wire id04471;
  wire id04472;
  wire id04473;
  wire id04474;
  wire id04475;
  wire id04476;
  wire id04477;
  wire id04478;
  wire id04479;
  wire id04480;
  wire id04481;
  wire id04482;
  wire id04483;
  wire id04484;
  wire id04485;
  wire id04486;
  wire id04487;
  wire id04488;
  wire id04489;
  wire id04490;
  wire id04491;
  wire id04492;
  wire id04493;
  wire id04494;
  wire id04495;
  wire id04496;
  wire id04497;
  wire id04498;
  wire id04499;
  wire id04500;
  wire id04501;
  wire id04502;
  wire id04503;
  wire id04504;
  wire id04505;
  wire id04506;
  wire id04507;
  wire id04508;
  wire id04509;
  wire id04510;
  wire id04511;
  wire id04512;
  wire id04513;
  wire id04514;
  wire id04515;
  wire id04516;
  wire id04517;
  wire id04518;
  wire id04519;
  wire id04520;
  wire id04521;
  wire id04522;
  wire id04523;
  wire id04524;
  wire id04525;
  wire id04526;
  wire id04527;
  wire id04528;
  wire id04529;
  wire id04530;
  wire id04531;
  wire id04532;
  wire id04533;
  wire id04534;
  wire id04535;
  wire id04536;
  wire id04537;
  wire id04538;
  wire id04539;
  wire id04540;
  wire id04541;
  wire id04542;
  wire id04543;
  wire id04544;
  wire id04545;
  wire id04546;
  wire id04547;
  wire id04548;
  wire id04549;
  wire id04550;
  wire id04551;
  wire id04552;
  wire id04553;
  wire id04554;
  wire id04555;
  wire id04556;
  wire id04557;
  wire id04558;
  wire id04559;
  wire id04560;
  wire id04561;
  wire id04562;
  wire id04563;
  wire id04564;
  wire id04565;
  wire id04566;
  wire id04567;
  wire id04568;
  wire id04569;
  wire id04570;
  wire id04571;
  wire id04572;
  wire id04573;
  wire id04574;
  wire id04575;
  wire id04576;
  wire id04577;
  wire id04578;
  wire id04579;
  wire id04580;
  wire id04581;
  wire id04582;
  wire id04583;
  wire id04584;
  wire id04585;
  wire id04586;
  wire id04587;
  wire id04588;
  wire id04589;
  wire id04590;
  wire id04591;
  wire id04592;
  wire id04593;
  wire id04594;
  wire id04595;
  wire id04596;
  wire id04597;
  wire id04598;
  wire id04599;
  wire id04600;
  wire id04601;
  wire id04602;
  wire id04603;
  wire id04604;
  wire id04605;
  wire id04606;
  wire id04607;
  wire id04608;
  wire id04609;
  wire id04610;
  wire id04611;
  wire id04612;
  wire id04613;
  wire id04614;
  wire id04615;
  wire id04616;
  wire id04617;
  wire id04618;
  wire id04619;
  wire id04620;
  wire id04621;
  wire id04622;
  wire id04623;
  wire id04624;
  wire id04625;
  wire id04626;
  wire id04627;
  wire id04628;
  wire id04629;
  wire id04630;
  wire id04631;
  wire id04632;
  wire id04633;
  wire id04634;
  wire id04635;
  wire id04636;
  wire id04637;
  wire id04638;
  wire id04639;
  wire id04640;
  wire id04641;
  wire id04642;
  wire id04643;
  wire id04644;
  wire id04645;
  wire id04646;
  wire id04647;
  wire id04648;
  wire id04649;
  wire id04650;
  wire id04651;
  wire id04652;
  wire id04653;
  wire id04654;
  wire id04655;
  wire id04656;
  wire id04657;
  wire id04658;
  wire id04659;
  wire id04660;
  wire id04661;
  wire id04662;
  wire id04663;
  wire id04664;
  wire id04665;
  wire id04666;
  wire id04667;
  wire id04668;
  wire id04669;
  wire id04670;
  wire id04671;
  wire id04672;
  wire id04673;
  wire id04674;
  wire id04675;
  wire id04676;
  wire id04677;
  wire id04678;
  wire id04679;
  wire id04680;
  wire id04681;
  wire id04682;
  wire id04683;
  wire id04684;
  wire id04685;
  wire id04686;
  wire id04687;
  wire id04688;
  wire id04689;
  wire id04690;
  wire id04691;
  wire id04692;
  wire id04693;
  wire id04694;
  wire id04695;
  wire id04696;
  wire id04697;
  wire id04698;
  wire id04699;
  wire id04700;
  wire id04701;
  wire id04702;
  wire id04703;
  wire id04704;
  wire id04705;
  wire id04706;
  wire id04707;
  wire id04708;
  wire id04709;
  wire id04710;
  wire id04711;
  wire id04712;
  wire id04713;
  wire id04714;
  wire id04715;
  wire id04716;
  wire id04717;
  wire id04718;
  wire id04719;
  wire id04720;
  wire id04721;
  wire id04722;
  wire id04723;
  wire id04724;
  wire id04725;
  wire id04726;
  wire id04727;
  wire id04728;
  wire id04729;
  wire id04730;
  wire id04731;
  wire id04732;
  wire id04733;
  wire id04734;
  wire id04735;
  wire id04736;
  wire id04737;
  wire id04738;
  wire id04739;
  wire id04740;
  wire id04741;
  wire id04742;
  wire id04743;
  wire id04744;
  wire id04745;
  wire id04746;
  wire id04747;
  wire id04748;
  wire id04749;
  wire id04750;
  wire id04751;
  wire id04752;
  wire id04753;
  wire id04754;
  wire id04755;
  wire id04756;
  wire id04757;
  wire id04758;
  wire id04759;
  wire id04760;
  wire id04761;
  wire id04762;
  wire id04763;
  wire id04764;
  wire id04765;
  wire id04766;
  wire id04767;
  wire id04768;
  wire id04769;
  wire id04770;
  wire id04771;
  wire id04772;
  wire id04773;
  wire id04774;
  wire id04775;
  wire id04776;
  wire id04777;
  wire id04778;
  wire id04779;
  wire id04780;
  wire id04781;
  wire id04782;
  wire id04783;
  wire id04784;
  wire id04785;
  wire id04786;
  wire id04787;
  wire id04788;
  wire id04789;
  wire id04790;
  wire id04791;
  wire id04792;
  wire id04793;
  wire id04794;
  wire id04795;
  wire id04796;
  wire id04797;
  wire id04798;
  wire id04799;
  wire id04800;
  wire id04801;
  wire id04802;
  wire id04803;
  wire id04804;
  wire id04805;
  wire id04806;
  wire id04807;
  wire id04808;
  wire id04809;
  wire id04810;
  wire id04811;
  wire id04812;
  wire id04813;
  wire id04814;
  wire id04815;
  wire id04816;
  wire id04817;
  wire id04818;
  wire id04819;
  wire id04820;
  wire id04821;
  wire id04822;
  wire id04823;
  wire id04824;
  wire id04825;
  wire id04826;
  wire id04827;
  wire id04828;
  wire id04829;
  wire id04830;
  wire id04831;
  wire id04832;
  wire id04833;
  wire id04834;
  wire id04835;
  wire id04836;
  wire id04837;
  wire id04838;
  wire id04839;
  wire id04840;
  wire id04841;
  wire id04842;
  wire id04843;
  wire id04844;
  wire id04845;
  wire id04846;
  wire id04847;
  wire id04848;
  wire id04849;
  wire id04850;
  wire id04851;
  wire id04852;
  wire id04853;
  wire id04854;
  wire id04855;
  wire id04856;
  wire id04857;
  wire id04858;
  wire \net_Buf-pad-result[1] ;
  wire \net_Buf-pad-result[0] ;
  wire \net_Buf-pad-result[3] ;
  wire \net_Buf-pad-result[2] ;


  defparam id00001.INIT = 8'hE8;
  LUT3 id00001 (
    .ADR0(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x2 ),
    .O(id04793)
  );

  defparam id00002.INIT = 16'h7117;
  LUT4 id00002 (
    .ADR0(id04775),
    .ADR1(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x0 ),
    .ADR2(id04770),
    .ADR3(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x3 ),
    .O(id04790)
  );

  defparam id00003.INIT = 16'h9669;
  LUT4 id00003 (
    .ADR0(id04794),
    .ADR1(id04791),
    .ADR2(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x3 ),
    .O(id04787)
  );

  defparam id00004.INIT = 4'h6;
  LUT2 id00004 (
    .ADR0(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x2 ),
    .O(id04794)
  );

  defparam id00005.INIT = 8'hE8;
  LUT3 id00005 (
    .ADR0(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x2 ),
    .O(id04791)
  );

  defparam id00006.INIT = 8'h71;
  LUT3 id00006 (
    .ADR0(id04834),
    .ADR1(id04832),
    .ADR2(id04831),
    .O(id04749)
  );

  defparam id00007.INIT = 8'hB2;
  LUT3 id00007 (
    .ADR0(id04850),
    .ADR1(id04847),
    .ADR2(id04848),
    .O(id04765)
  );

  defparam id00008.INIT = 16'hE817;
  LUT4 id00008 (
    .ADR0(id04776),
    .ADR1(id04764),
    .ADR2(id04761),
    .ADR3(id04792),
    .O(\net_Buf-pad-result[33] )
  );

  defparam id00009.INIT = 4'h9;
  LUT2 id00009 (
    .ADR0(id04783),
    .ADR1(id04784),
    .O(id04792)
  );

  defparam id00010.INIT = 4'h4;
  LUT2 id00010 (
    .ADR0(id04762),
    .ADR1(id04767),
    .O(id04783)
  );

  defparam id00011.INIT = 4'h9;
  LUT2 id00011 (
    .ADR0(id04781),
    .ADR1(id04782),
    .O(id04784)
  );

  defparam id00012.INIT = 8'h3A;
  LUT3 id00012 (
    .ADR0(id04765),
    .ADR1(id04753),
    .ADR2(id04768),
    .O(id04781)
  );

  defparam id00013.INIT = 4'h6;
  LUT2 id00013 (
    .ADR0(id04785),
    .ADR1(id04786),
    .O(id04782)
  );

  defparam id00014.INIT = 16'h9669;
  LUT4 id00014 (
    .ADR0(id03658),
    .ADR1(id04779),
    .ADR2(id04778),
    .ADR3(id04777),
    .O(id04785)
  );

  defparam id00015.INIT = 8'hC5;
  LUT3 id00015 (
    .ADR0(id04747),
    .ADR1(id04759),
    .ADR2(id04754),
    .O(id03658)
  );

  defparam id00016.INIT = 4'h6;
  LUT2 id00016 (
    .ADR0(id04780),
    .ADR1(id03577),
    .O(id04779)
  );

  defparam id00017.INIT = 16'h6996;
  LUT4 id00017 (
    .ADR0(id03576),
    .ADR1(id03571),
    .ADR2(id03570),
    .ADR3(id03573),
    .O(id04780)
  );

  defparam id00018.INIT = 8'h35;
  LUT3 id00018 (
    .ADR0(id04745),
    .ADR1(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x0 ),
    .ADR2(id04748),
    .O(id03576)
  );

  defparam id00019.INIT = 4'h9;
  LUT2 id00019 (
    .ADR0(id03572),
    .ADR1(id03453),
    .O(id03571)
  );

  defparam id00020.INIT = 16'h9669;
  LUT4 id00020 (
    .ADR0(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x2 ),
    .O(id03572)
  );

  defparam id00021.INIT = 8'hE8;
  LUT3 id00021 (
    .ADR0(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x2 ),
    .O(id03453)
  );

  defparam id00022.INIT = 16'h7117;
  LUT4 id00022 (
    .ADR0(id04751),
    .ADR1(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x0 ),
    .ADR2(id04746),
    .ADR3(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x3 ),
    .O(id03570)
  );

  defparam id00023.INIT = 16'h6996;
  LUT4 id00023 (
    .ADR0(id03452),
    .ADR1(id03455),
    .ADR2(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x3 ),
    .O(id03573)
  );

  defparam id00024.INIT = 4'h6;
  LUT2 id00024 (
    .ADR0(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x2 ),
    .O(id03452)
  );

  defparam id00025.INIT = 8'hE8;
  LUT3 id00025 (
    .ADR0(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x2 ),
    .O(id03455)
  );

  defparam id00026.INIT = 8'h71;
  LUT3 id00026 (
    .ADR0(id04760),
    .ADR1(id04758),
    .ADR2(id04757),
    .O(id03577)
  );

  defparam id00027.INIT = 8'h3A;
  LUT3 id00027 (
    .ADR0(id04787),
    .ADR1(id04749),
    .ADR2(id04752),
    .O(id04778)
  );

  defparam id00028.INIT = 4'h9;
  LUT2 id00028 (
    .ADR0(id03454),
    .ADR1(id03449),
    .O(id04777)
  );

  defparam id00029.INIT = 16'h9669;
  LUT4 id00029 (
    .ADR0(id03448),
    .ADR1(id03451),
    .ADR2(id03450),
    .ADR3(id03461),
    .O(id03454)
  );

  defparam id00030.INIT = 8'h35;
  LUT3 id00030 (
    .ADR0(id04793),
    .ADR1(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x0 ),
    .ADR2(id04788),
    .O(id03448)
  );

  defparam id00031.INIT = 4'h9;
  LUT2 id00031 (
    .ADR0(id03460),
    .ADR1(id03463),
    .O(id03451)
  );

  defparam id00032.INIT = 16'h9669;
  LUT4 id00032 (
    .ADR0(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x2 ),
    .O(id03460)
  );

  defparam id00033.INIT = 8'hE8;
  LUT3 id00033 (
    .ADR0(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x2 ),
    .O(id03463)
  );

  defparam id00034.INIT = 16'h8EE8;
  LUT4 id00034 (
    .ADR0(id04791),
    .ADR1(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .ADR2(id04794),
    .ADR3(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x3 ),
    .O(id03450)
  );

  defparam id00035.INIT = 16'h9669;
  LUT4 id00035 (
    .ADR0(id03462),
    .ADR1(id03457),
    .ADR2(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x3 ),
    .O(id03461)
  );

  defparam id00036.INIT = 4'h6;
  LUT2 id00036 (
    .ADR0(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x2 ),
    .O(id03462)
  );

  defparam id00037.INIT = 8'hE8;
  LUT3 id00037 (
    .ADR0(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x2 ),
    .O(id03457)
  );

  defparam id00038.INIT = 8'h71;
  LUT3 id00038 (
    .ADR0(id04750),
    .ADR1(id04790),
    .ADR2(id04789),
    .O(id03449)
  );

  defparam id00039.INIT = 8'hB2;
  LUT3 id00039 (
    .ADR0(id04766),
    .ADR1(id04755),
    .ADR2(id04756),
    .O(id04786)
  );

  defparam id00040.INIT = 4'h9;
  LUT2 id00040 (
    .ADR0(id03456),
    .ADR1(id03459),
    .O(\net_Buf-pad-result[34] )
  );

  defparam id00041.INIT = 16'h00BF;
  LUT4 id00041 (
    .ADR0(id04792),
    .ADR1(id04773),
    .ADR2(id04776),
    .ADR3(id03458),
    .O(id03456)
  );

  defparam id00042.INIT = 16'hB200;
  LUT4 id00042 (
    .ADR0(id04764),
    .ADR1(id04762),
    .ADR2(id04767),
    .ADR3(id04784),
    .O(id03458)
  );

  defparam id00043.INIT = 4'h6;
  LUT2 id00043 (
    .ADR0(id03469),
    .ADR1(id03180),
    .O(id03459)
  );

  defparam id00044.INIT = 4'h4;
  LUT2 id00044 (
    .ADR0(id04781),
    .ADR1(id04782),
    .O(id03469)
  );

  defparam id00045.INIT = 4'h9;
  LUT2 id00045 (
    .ADR0(id03167),
    .ADR1(id03173),
    .O(id03180)
  );

  defparam id00046.INIT = 8'h3A;
  LUT3 id00046 (
    .ADR0(id04786),
    .ADR1(id04777),
    .ADR2(id04785),
    .O(id03167)
  );

  defparam id00047.INIT = 4'h6;
  LUT2 id00047 (
    .ADR0(id03162),
    .ADR1(id03165),
    .O(id03173)
  );

  defparam id00048.INIT = 16'h9669;
  LUT4 id00048 (
    .ADR0(id03164),
    .ADR1(id03174),
    .ADR2(id03176),
    .ADR3(id03175),
    .O(id03162)
  );

  defparam id00049.INIT = 8'h35;
  LUT3 id00049 (
    .ADR0(id03573),
    .ADR1(id03577),
    .ADR2(id04780),
    .O(id03164)
  );

  defparam id00050.INIT = 4'h9;
  LUT2 id00050 (
    .ADR0(id03170),
    .ADR1(id03169),
    .O(id03174)
  );

  defparam id00051.INIT = 16'h6996;
  LUT4 id00051 (
    .ADR0(id03172),
    .ADR1(id03171),
    .ADR2(id03219),
    .ADR3(id03218),
    .O(id03170)
  );

  defparam id00052.INIT = 8'h35;
  LUT3 id00052 (
    .ADR0(id03453),
    .ADR1(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x0 ),
    .ADR2(id03572),
    .O(id03172)
  );

  defparam id00053.INIT = 4'h9;
  LUT2 id00053 (
    .ADR0(id03221),
    .ADR1(id03220),
    .O(id03171)
  );

  defparam id00054.INIT = 16'h9669;
  LUT4 id00054 (
    .ADR0(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x2 ),
    .O(id03221)
  );

  defparam id00055.INIT = 8'hE8;
  LUT3 id00055 (
    .ADR0(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x2 ),
    .O(id03220)
  );

  defparam id00056.INIT = 16'h7117;
  LUT4 id00056 (
    .ADR0(id03455),
    .ADR1(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x0 ),
    .ADR2(id03452),
    .ADR3(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x3 ),
    .O(id03219)
  );

  defparam id00057.INIT = 16'h6996;
  LUT4 id00057 (
    .ADR0(id03215),
    .ADR1(id03214),
    .ADR2(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x3 ),
    .O(id03218)
  );

  defparam id00058.INIT = 4'h6;
  LUT2 id00058 (
    .ADR0(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x2 ),
    .O(id03215)
  );

  defparam id00059.INIT = 8'hE8;
  LUT3 id00059 (
    .ADR0(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x2 ),
    .O(id03214)
  );

  defparam id00060.INIT = 8'hB2;
  LUT3 id00060 (
    .ADR0(id03576),
    .ADR1(id03571),
    .ADR2(id03570),
    .O(id03169)
  );

  defparam id00061.INIT = 8'hC5;
  LUT3 id00061 (
    .ADR0(id03449),
    .ADR1(id03461),
    .ADR2(id03454),
    .O(id03176)
  );

  defparam id00062.INIT = 4'h6;
  LUT2 id00062 (
    .ADR0(id03217),
    .ADR1(id03216),
    .O(id03175)
  );

  defparam id00063.INIT = 16'h9669;
  LUT4 id00063 (
    .ADR0(id03227),
    .ADR1(id03226),
    .ADR2(id03229),
    .ADR3(id03228),
    .O(id03217)
  );

  defparam id00064.INIT = 8'h35;
  LUT3 id00064 (
    .ADR0(id03463),
    .ADR1(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x0 ),
    .ADR2(id03460),
    .O(id03227)
  );

  defparam id00065.INIT = 4'h9;
  LUT2 id00065 (
    .ADR0(id03223),
    .ADR1(id03222),
    .O(id03226)
  );

  defparam id00066.INIT = 16'h9669;
  LUT4 id00066 (
    .ADR0(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x2 ),
    .O(id03223)
  );

  defparam id00067.INIT = 8'hE8;
  LUT3 id00067 (
    .ADR0(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x2 ),
    .O(id03222)
  );

  defparam id00068.INIT = 16'h8EE8;
  LUT4 id00068 (
    .ADR0(id03457),
    .ADR1(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .ADR2(id03462),
    .ADR3(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x3 ),
    .O(id03229)
  );

  defparam id00069.INIT = 16'h6996;
  LUT4 id00069 (
    .ADR0(id03225),
    .ADR1(id03224),
    .ADR2(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x3 ),
    .O(id03228)
  );

  defparam id00070.INIT = 4'h6;
  LUT2 id00070 (
    .ADR0(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x2 ),
    .O(id03225)
  );

  defparam id00071.INIT = 8'hE8;
  LUT3 id00071 (
    .ADR0(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x2 ),
    .O(id03224)
  );

  defparam id00072.INIT = 8'hD4;
  LUT3 id00072 (
    .ADR0(id03448),
    .ADR1(id03451),
    .ADR2(id03450),
    .O(id03216)
  );

  defparam id00073.INIT = 8'hB2;
  LUT3 id00073 (
    .ADR0(id03658),
    .ADR1(id04779),
    .ADR2(id04778),
    .O(id03165)
  );

  defparam id00074.INIT = 16'h2BD4;
  LUT4 id00074 (
    .ADR0(id03456),
    .ADR1(id03469),
    .ADR2(id03180),
    .ADR3(id03235),
    .O(\net_Buf-pad-result[35] )
  );

  defparam id00075.INIT = 4'h6;
  LUT2 id00075 (
    .ADR0(id03234),
    .ADR1(id03237),
    .O(id03235)
  );

  defparam id00076.INIT = 4'h4;
  LUT2 id00076 (
    .ADR0(id03167),
    .ADR1(id03173),
    .O(id03234)
  );

  defparam id00077.INIT = 4'h9;
  LUT2 id00077 (
    .ADR0(id03592),
    .ADR1(id03587),
    .O(id03237)
  );

  defparam id00078.INIT = 8'h3A;
  LUT3 id00078 (
    .ADR0(id03165),
    .ADR1(id03175),
    .ADR2(id03162),
    .O(id03592)
  );

  defparam id00079.INIT = 4'h6;
  LUT2 id00079 (
    .ADR0(id03595),
    .ADR1(id03594),
    .O(id03587)
  );

  defparam id00080.INIT = 16'h9669;
  LUT4 id00080 (
    .ADR0(id03588),
    .ADR1(id03599),
    .ADR2(id03598),
    .ADR3(id03600),
    .O(id03595)
  );

  defparam id00081.INIT = 8'hC5;
  LUT3 id00081 (
    .ADR0(id03218),
    .ADR1(id03169),
    .ADR2(id03170),
    .O(id03588)
  );

  defparam id00082.INIT = 4'h6;
  LUT2 id00082 (
    .ADR0(id03597),
    .ADR1(id03596),
    .O(id03599)
  );

  defparam id00083.INIT = 16'h6996;
  LUT4 id00083 (
    .ADR0(id03606),
    .ADR1(id03605),
    .ADR2(id03608),
    .ADR3(id03607),
    .O(id03597)
  );

  defparam id00084.INIT = 8'h35;
  LUT3 id00084 (
    .ADR0(id03220),
    .ADR1(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x0 ),
    .ADR2(id03221),
    .O(id03606)
  );

  defparam id00085.INIT = 4'h9;
  LUT2 id00085 (
    .ADR0(id03602),
    .ADR1(id03601),
    .O(id03605)
  );

  defparam id00086.INIT = 16'h9669;
  LUT4 id00086 (
    .ADR0(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x2 ),
    .O(id03602)
  );

  defparam id00087.INIT = 8'hE8;
  LUT3 id00087 (
    .ADR0(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x2 ),
    .O(id03601)
  );

  defparam id00088.INIT = 16'h7117;
  LUT4 id00088 (
    .ADR0(id03214),
    .ADR1(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x0 ),
    .ADR2(id03215),
    .ADR3(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x3 ),
    .O(id03608)
  );

  defparam id00089.INIT = 16'h6996;
  LUT4 id00089 (
    .ADR0(id03604),
    .ADR1(id03603),
    .ADR2(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x3 ),
    .O(id03607)
  );

  defparam id00090.INIT = 4'h6;
  LUT2 id00090 (
    .ADR0(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x2 ),
    .O(id03604)
  );

  defparam id00091.INIT = 8'hE8;
  LUT3 id00091 (
    .ADR0(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x2 ),
    .O(id03603)
  );

  defparam id00092.INIT = 8'h71;
  LUT3 id00092 (
    .ADR0(id03172),
    .ADR1(id03219),
    .ADR2(id03171),
    .O(id03596)
  );

  defparam id00093.INIT = 8'h35;
  LUT3 id00093 (
    .ADR0(id03228),
    .ADR1(id03216),
    .ADR2(id03217),
    .O(id03598)
  );

  defparam id00094.INIT = 4'h9;
  LUT2 id00094 (
    .ADR0(id03551),
    .ADR1(id03550),
    .O(id03600)
  );

  defparam id00095.INIT = 16'h9669;
  LUT4 id00095 (
    .ADR0(id03553),
    .ADR1(id03552),
    .ADR2(id03547),
    .ADR3(id03546),
    .O(id03551)
  );

  defparam id00096.INIT = 8'h35;
  LUT3 id00096 (
    .ADR0(id03222),
    .ADR1(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x0 ),
    .ADR2(id03223),
    .O(id03553)
  );

  defparam id00097.INIT = 4'h9;
  LUT2 id00097 (
    .ADR0(id03549),
    .ADR1(id03548),
    .O(id03552)
  );

  defparam id00098.INIT = 16'h9669;
  LUT4 id00098 (
    .ADR0(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x2 ),
    .O(id03549)
  );

  defparam id00099.INIT = 8'hE8;
  LUT3 id00099 (
    .ADR0(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x2 ),
    .O(id03548)
  );

  defparam id00100.INIT = 16'h7117;
  LUT4 id00100 (
    .ADR0(id03224),
    .ADR1(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x0 ),
    .ADR2(id03225),
    .ADR3(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x3 ),
    .O(id03547)
  );

  defparam id00101.INIT = 16'h6996;
  LUT4 id00101 (
    .ADR0(id03559),
    .ADR1(id03558),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x3 ),
    .O(id03546)
  );

  defparam id00102.INIT = 4'h6;
  LUT2 id00102 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x2 ),
    .O(id03559)
  );

  defparam id00103.INIT = 8'hE8;
  LUT3 id00103 (
    .ADR0(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x2 ),
    .O(id03558)
  );

  defparam id00104.INIT = 8'hD4;
  LUT3 id00104 (
    .ADR0(id03227),
    .ADR1(id03226),
    .ADR2(id03229),
    .O(id03550)
  );

  defparam id00105.INIT = 8'hB2;
  LUT3 id00105 (
    .ADR0(id03164),
    .ADR1(id03174),
    .ADR2(id03176),
    .O(id03594)
  );

  defparam id00106.INIT = 4'h9;
  LUT2 id00106 (
    .ADR0(id03561),
    .ADR1(id03560),
    .O(\net_Buf-pad-result[36] )
  );

  defparam id00107.INIT = 16'hBF00;
  LUT4 id00107 (
    .ADR0(id03456),
    .ADR1(id03235),
    .ADR2(id03459),
    .ADR3(id03555),
    .O(id03561)
  );

  defparam id00108.INIT = 16'h07FF;
  LUT4 id00108 (
    .ADR0(id03469),
    .ADR1(id03180),
    .ADR2(id03234),
    .ADR3(id03237),
    .O(id03555)
  );

  defparam id00109.INIT = 4'h6;
  LUT2 id00109 (
    .ADR0(id03554),
    .ADR1(id03557),
    .O(id03560)
  );

  defparam id00110.INIT = 4'h4;
  LUT2 id00110 (
    .ADR0(id03592),
    .ADR1(id03587),
    .O(id03554)
  );

  defparam id00111.INIT = 4'h9;
  LUT2 id00111 (
    .ADR0(id03494),
    .ADR1(id03520),
    .O(id03557)
  );

  defparam id00112.INIT = 8'h3A;
  LUT3 id00112 (
    .ADR0(id03594),
    .ADR1(id03600),
    .ADR2(id03595),
    .O(id03494)
  );

  defparam id00113.INIT = 4'h9;
  LUT2 id00113 (
    .ADR0(id03495),
    .ADR1(id03499),
    .O(id03520)
  );

  defparam id00114.INIT = 16'h6996;
  LUT4 id00114 (
    .ADR0(id03501),
    .ADR1(id03491),
    .ADR2(id03513),
    .ADR3(id03507),
    .O(id03495)
  );

  defparam id00115.INIT = 8'h35;
  LUT3 id00115 (
    .ADR0(id03607),
    .ADR1(id03596),
    .ADR2(id03597),
    .O(id03501)
  );

  defparam id00116.INIT = 4'h9;
  LUT2 id00116 (
    .ADR0(id03509),
    .ADR1(id03583),
    .O(id03491)
  );

  defparam id00117.INIT = 16'h6996;
  LUT4 id00117 (
    .ADR0(id03585),
    .ADR1(id03579),
    .ADR2(id03581),
    .ADR3(id03591),
    .O(id03509)
  );

  defparam id00118.INIT = 8'h35;
  LUT3 id00118 (
    .ADR0(id03601),
    .ADR1(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x0 ),
    .ADR2(id03602),
    .O(id03585)
  );

  defparam id00119.INIT = 4'h9;
  LUT2 id00119 (
    .ADR0(id03504),
    .ADR1(id03464),
    .O(id03579)
  );

  defparam id00120.INIT = 16'h9669;
  LUT4 id00120 (
    .ADR0(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x2 ),
    .O(id03504)
  );

  defparam id00121.INIT = 8'hE8;
  LUT3 id00121 (
    .ADR0(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x2 ),
    .O(id03464)
  );

  defparam id00122.INIT = 16'h7117;
  LUT4 id00122 (
    .ADR0(id03603),
    .ADR1(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x0 ),
    .ADR2(id03604),
    .ADR3(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x3 ),
    .O(id03581)
  );

  defparam id00123.INIT = 16'h6996;
  LUT4 id00123 (
    .ADR0(id03473),
    .ADR1(id03255),
    .ADR2(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x3 ),
    .O(id03591)
  );

  defparam id00124.INIT = 4'h6;
  LUT2 id00124 (
    .ADR0(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x2 ),
    .O(id03473)
  );

  defparam id00125.INIT = 8'hE8;
  LUT3 id00125 (
    .ADR0(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x2 ),
    .O(id03255)
  );

  defparam id00126.INIT = 8'hB2;
  LUT3 id00126 (
    .ADR0(id03606),
    .ADR1(id03605),
    .ADR2(id03608),
    .O(id03583)
  );

  defparam id00127.INIT = 8'h35;
  LUT3 id00127 (
    .ADR0(id03550),
    .ADR1(id03546),
    .ADR2(id03551),
    .O(id03513)
  );

  defparam id00128.INIT = 4'h9;
  LUT2 id00128 (
    .ADR0(id03470),
    .ADR1(id03472),
    .O(id03507)
  );

  defparam id00129.INIT = 16'h9669;
  LUT4 id00129 (
    .ADR0(id03420),
    .ADR1(id03423),
    .ADR2(id03417),
    .ADR3(id03419),
    .O(id03470)
  );

  defparam id00130.INIT = 8'h35;
  LUT3 id00130 (
    .ADR0(id03548),
    .ADR1(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x0 ),
    .ADR2(id03549),
    .O(id03420)
  );

  defparam id00131.INIT = 4'h9;
  LUT2 id00131 (
    .ADR0(id03429),
    .ADR1(id03475),
    .O(id03423)
  );

  defparam id00132.INIT = 16'h9669;
  LUT4 id00132 (
    .ADR0(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x2 ),
    .O(id03429)
  );

  defparam id00133.INIT = 8'hE8;
  LUT3 id00133 (
    .ADR0(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x2 ),
    .O(id03475)
  );

  defparam id00134.INIT = 16'h7117;
  LUT4 id00134 (
    .ADR0(id03558),
    .ADR1(GND_NET),
    .ADR2(id03559),
    .ADR3(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x3 ),
    .O(id03417)
  );

  defparam id00135.INIT = 8'h96;
  LUT3 id00135 (
    .ADR0(id03430),
    .ADR1(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 ),
    .O(id03419)
  );

  defparam id00136.INIT = 8'hE8;
  LUT3 id00136 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x2 ),
    .O(id03430)
  );

  defparam id00137.INIT = 8'h71;
  LUT3 id00137 (
    .ADR0(id03553),
    .ADR1(id03547),
    .ADR2(id03552),
    .O(id03472)
  );

  defparam id00138.INIT = 8'hB2;
  LUT3 id00138 (
    .ADR0(id03588),
    .ADR1(id03599),
    .ADR2(id03598),
    .O(id03499)
  );

  defparam id00139.INIT = 16'h0BF4;
  LUT4 id00139 (
    .ADR0(id03561),
    .ADR1(id03560),
    .ADR2(id03424),
    .ADR3(id03426),
    .O(\net_Buf-pad-result[37] )
  );

  defparam id00140.INIT = 4'h6;
  LUT2 id00140 (
    .ADR0(id03436),
    .ADR1(id03438),
    .O(id03426)
  );

  defparam id00141.INIT = 4'h9;
  LUT2 id00141 (
    .ADR0(id03432),
    .ADR1(id03434),
    .O(id03436)
  );

  defparam id00142.INIT = 4'h9;
  LUT2 id00142 (
    .ADR0(id03444),
    .ADR1(id03446),
    .O(id03432)
  );

  defparam id00143.INIT = 16'h6996;
  LUT4 id00143 (
    .ADR0(id03440),
    .ADR1(id03442),
    .ADR2(id03479),
    .ADR3(id03481),
    .O(id03444)
  );

  defparam id00144.INIT = 4'h9;
  LUT2 id00144 (
    .ADR0(id03257),
    .ADR1(id03256),
    .O(id03440)
  );

  defparam id00145.INIT = 8'h69;
  LUT3 id00145 (
    .ADR0(id03259),
    .ADR1(id03258),
    .ADR2(id03260),
    .O(id03257)
  );

  defparam id00146.INIT = 4'h6;
  LUT2 id00146 (
    .ADR0(id03497),
    .ADR1(id03492),
    .O(id03259)
  );

  defparam id00147.INIT = 8'h60;
  LUT3 id00147 (
    .ADR0(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 ),
    .ADR2(id03430),
    .O(id03492)
  );

  defparam id00148.INIT = 16'h8778;
  LUT4 id00148 (
    .ADR0(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 ),
    .ADR2(\u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 ),
    .ADR3(VCC_NET),
    .O(id03497)
  );

  defparam id00149.INIT = 8'h35;
  LUT3 id00149 (
    .ADR0(id03475),
    .ADR1(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x0 ),
    .ADR2(id03429),
    .O(id03258)
  );

  defparam id00150.INIT = 4'h9;
  LUT2 id00150 (
    .ADR0(id03493),
    .ADR1(id03496),
    .O(id03260)
  );

  defparam id00151.INIT = 16'h9669;
  LUT4 id00151 (
    .ADR0(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x2 ),
    .O(id03493)
  );

  defparam id00152.INIT = 8'hE8;
  LUT3 id00152 (
    .ADR0(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x2 ),
    .O(id03496)
  );

  defparam id00153.INIT = 8'hB2;
  LUT3 id00153 (
    .ADR0(id03420),
    .ADR1(id03423),
    .ADR2(id03417),
    .O(id03256)
  );

  defparam id00154.INIT = 8'hC5;
  LUT3 id00154 (
    .ADR0(id03591),
    .ADR1(id03583),
    .ADR2(id03509),
    .O(id03442)
  );

  defparam id00155.INIT = 4'h9;
  LUT2 id00155 (
    .ADR0(id03498),
    .ADR1(id03503),
    .O(id03479)
  );

  defparam id00156.INIT = 16'h6996;
  LUT4 id00156 (
    .ADR0(id03500),
    .ADR1(id03502),
    .ADR2(id03511),
    .ADR3(id03510),
    .O(id03498)
  );

  defparam id00157.INIT = 8'h35;
  LUT3 id00157 (
    .ADR0(id03464),
    .ADR1(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x0 ),
    .ADR2(id03504),
    .O(id03500)
  );

  defparam id00158.INIT = 4'h9;
  LUT2 id00158 (
    .ADR0(id03505),
    .ADR1(id03512),
    .O(id03502)
  );

  defparam id00159.INIT = 16'h9669;
  LUT4 id00159 (
    .ADR0(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x2 ),
    .O(id03505)
  );

  defparam id00160.INIT = 8'hE8;
  LUT3 id00160 (
    .ADR0(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x2 ),
    .O(id03512)
  );

  defparam id00161.INIT = 16'h7117;
  LUT4 id00161 (
    .ADR0(id03255),
    .ADR1(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x0 ),
    .ADR2(id03473),
    .ADR3(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x3 ),
    .O(id03511)
  );

  defparam id00162.INIT = 16'h6996;
  LUT4 id00162 (
    .ADR0(id03506),
    .ADR1(id03508),
    .ADR2(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x3 ),
    .O(id03510)
  );

  defparam id00163.INIT = 4'h6;
  LUT2 id00163 (
    .ADR0(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x2 ),
    .O(id03506)
  );

  defparam id00164.INIT = 8'hE8;
  LUT3 id00164 (
    .ADR0(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x2 ),
    .O(id03508)
  );

  defparam id00165.INIT = 8'hB2;
  LUT3 id00165 (
    .ADR0(id03585),
    .ADR1(id03579),
    .ADR2(id03581),
    .O(id03503)
  );

  defparam id00166.INIT = 8'h35;
  LUT3 id00166 (
    .ADR0(id03472),
    .ADR1(id03419),
    .ADR2(id03470),
    .O(id03481)
  );

  defparam id00167.INIT = 8'hB2;
  LUT3 id00167 (
    .ADR0(id03501),
    .ADR1(id03491),
    .ADR2(id03513),
    .O(id03446)
  );

  defparam id00168.INIT = 8'hC5;
  LUT3 id00168 (
    .ADR0(id03507),
    .ADR1(id03499),
    .ADR2(id03495),
    .O(id03434)
  );

  defparam id00169.INIT = 4'h4;
  LUT2 id00169 (
    .ADR0(id03494),
    .ADR1(id03520),
    .O(id03438)
  );

  defparam id00170.INIT = 4'h8;
  LUT2 id00170 (
    .ADR0(id03554),
    .ADR1(id03557),
    .O(id03424)
  );

  defparam id00171.INIT = 8'h69;
  LUT3 id00171 (
    .ADR0(id03582),
    .ADR1(id03584),
    .ADR2(id03578),
    .O(\net_Buf-pad-result[38] )
  );

  defparam id00172.INIT = 16'hBF00;
  LUT4 id00172 (
    .ADR0(id03561),
    .ADR1(id03426),
    .ADR2(id03560),
    .ADR3(id03580),
    .O(id03582)
  );

  defparam id00173.INIT = 8'h1F;
  LUT3 id00173 (
    .ADR0(id03424),
    .ADR1(id03438),
    .ADR2(id03436),
    .O(id03580)
  );

  defparam id00174.INIT = 4'h4;
  LUT2 id00174 (
    .ADR0(id03434),
    .ADR1(id03432),
    .O(id03584)
  );

  defparam id00175.INIT = 4'h9;
  LUT2 id00175 (
    .ADR0(id03590),
    .ADR1(id03593),
    .O(id03578)
  );

  defparam id00176.INIT = 8'hC5;
  LUT3 id00176 (
    .ADR0(id03440),
    .ADR1(id03446),
    .ADR2(id03444),
    .O(id03590)
  );

  defparam id00177.INIT = 4'h6;
  LUT2 id00177 (
    .ADR0(id03467),
    .ADR1(id03465),
    .O(id03593)
  );

  defparam id00178.INIT = 16'h1EE1;
  LUT4 id00178 (
    .ADR0(id03468),
    .ADR1(id03246),
    .ADR2(id03586),
    .ADR3(id03478),
    .O(id03467)
  );

  defparam id00179.INIT = 4'h4;
  LUT2 id00179 (
    .ADR0(id03474),
    .ADR1(id03421),
    .O(id03468)
  );

  defparam id00180.INIT = 8'hC5;
  LUT3 id00180 (
    .ADR0(id03510),
    .ADR1(id03503),
    .ADR2(id03498),
    .O(id03474)
  );

  defparam id00181.INIT = 4'h6;
  LUT2 id00181 (
    .ADR0(id03422),
    .ADR1(id03416),
    .O(id03421)
  );

  defparam id00182.INIT = 16'h6996;
  LUT4 id00182 (
    .ADR0(id03418),
    .ADR1(id03428),
    .ADR2(id03431),
    .ADR3(id03425),
    .O(id03422)
  );

  defparam id00183.INIT = 8'h35;
  LUT3 id00183 (
    .ADR0(id03512),
    .ADR1(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x0 ),
    .ADR2(id03505),
    .O(id03418)
  );

  defparam id00184.INIT = 4'h9;
  LUT2 id00184 (
    .ADR0(id03427),
    .ADR1(id03437),
    .O(id03428)
  );

  defparam id00185.INIT = 16'h9669;
  LUT4 id00185 (
    .ADR0(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x2 ),
    .O(id03427)
  );

  defparam id00186.INIT = 8'hE8;
  LUT3 id00186 (
    .ADR0(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x2 ),
    .O(id03437)
  );

  defparam id00187.INIT = 16'h7117;
  LUT4 id00187 (
    .ADR0(id03508),
    .ADR1(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x0 ),
    .ADR2(id03506),
    .ADR3(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x3 ),
    .O(id03431)
  );

  defparam id00188.INIT = 16'h6996;
  LUT4 id00188 (
    .ADR0(id03439),
    .ADR1(id03433),
    .ADR2(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x3 ),
    .O(id03425)
  );

  defparam id00189.INIT = 4'h6;
  LUT2 id00189 (
    .ADR0(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x2 ),
    .O(id03439)
  );

  defparam id00190.INIT = 8'hE8;
  LUT3 id00190 (
    .ADR0(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x2 ),
    .O(id03433)
  );

  defparam id00191.INIT = 8'h71;
  LUT3 id00191 (
    .ADR0(id03500),
    .ADR1(id03511),
    .ADR2(id03502),
    .O(id03416)
  );

  defparam id00192.INIT = 4'h4;
  LUT2 id00192 (
    .ADR0(id03421),
    .ADR1(id03474),
    .O(id03246)
  );

  defparam id00193.INIT = 8'hC5;
  LUT3 id00193 (
    .ADR0(id03497),
    .ADR1(id03256),
    .ADR2(id03257),
    .O(id03586)
  );

  defparam id00194.INIT = 4'h6;
  LUT2 id00194 (
    .ADR0(id03435),
    .ADR1(id03445),
    .O(id03478)
  );

  defparam id00195.INIT = 16'h9669;
  LUT4 id00195 (
    .ADR0(id03447),
    .ADR1(id03441),
    .ADR2(id03443),
    .ADR3(id03480),
    .O(id03435)
  );

  defparam id00196.INIT = 8'h35;
  LUT3 id00196 (
    .ADR0(id03496),
    .ADR1(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x0 ),
    .ADR2(id03493),
    .O(id03447)
  );

  defparam id00197.INIT = 4'h9;
  LUT2 id00197 (
    .ADR0(id03482),
    .ADR1(id03517),
    .O(id03441)
  );

  defparam id00198.INIT = 16'h9669;
  LUT4 id00198 (
    .ADR0(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x2 ),
    .O(id03482)
  );

  defparam id00199.INIT = 8'hE8;
  LUT3 id00199 (
    .ADR0(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x2 ),
    .O(id03517)
  );

  defparam id00200.INIT = 16'h6000;
  LUT4 id00200 (
    .ADR0(\u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 ),
    .O(id03443)
  );

  defparam id00201.INIT = 8'h78;
  LUT3 id00201 (
    .ADR0(\u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[38].u_compressor42_cell.x3 ),
    .O(id03480)
  );

  defparam id00202.INIT = 8'hB2;
  LUT3 id00202 (
    .ADR0(id03492),
    .ADR1(id03258),
    .ADR2(id03260),
    .O(id03445)
  );

  defparam id00203.INIT = 8'hB2;
  LUT3 id00203 (
    .ADR0(id03442),
    .ADR1(id03479),
    .ADR2(id03481),
    .O(id03465)
  );

  defparam id00204.INIT = 8'h1E;
  LUT3 id00204 (
    .ADR0(id03527),
    .ADR1(id03187),
    .ADR2(id03515),
    .O(\net_Buf-pad-result[39] )
  );

  defparam id00205.INIT = 8'h2B;
  LUT3 id00205 (
    .ADR0(id03582),
    .ADR1(id03584),
    .ADR2(id03578),
    .O(id03515)
  );

  defparam id00206.INIT = 4'h8;
  LUT2 id00206 (
    .ADR0(id03529),
    .ADR1(id03523),
    .O(id03527)
  );

  defparam id00207.INIT = 4'h4;
  LUT2 id00207 (
    .ADR0(id03590),
    .ADR1(id03593),
    .O(id03529)
  );

  defparam id00208.INIT = 4'h9;
  LUT2 id00208 (
    .ADR0(id03525),
    .ADR1(id03535),
    .O(id03523)
  );

  defparam id00209.INIT = 8'h3A;
  LUT3 id00209 (
    .ADR0(id03465),
    .ADR1(id03478),
    .ADR2(id03467),
    .O(id03525)
  );

  defparam id00210.INIT = 4'h9;
  LUT2 id00210 (
    .ADR0(id03537),
    .ADR1(id03531),
    .O(id03535)
  );

  defparam id00211.INIT = 8'h0E;
  LUT3 id00211 (
    .ADR0(id03586),
    .ADR1(id03246),
    .ADR2(id03468),
    .O(id03537)
  );

  defparam id00212.INIT = 16'h6996;
  LUT4 id00212 (
    .ADR0(id03533),
    .ADR1(id03543),
    .ADR2(id03545),
    .ADR3(id03539),
    .O(id03531)
  );

  defparam id00213.INIT = 8'h35;
  LUT3 id00213 (
    .ADR0(id03425),
    .ADR1(id03416),
    .ADR2(id03422),
    .O(id03533)
  );

  defparam id00214.INIT = 4'h9;
  LUT2 id00214 (
    .ADR0(id03541),
    .ADR1(id03488),
    .O(id03543)
  );

  defparam id00215.INIT = 16'h6996;
  LUT4 id00215 (
    .ADR0(id03490),
    .ADR1(id03484),
    .ADR2(id03486),
    .ADR3(id03516),
    .O(id03541)
  );

  defparam id00216.INIT = 8'h35;
  LUT3 id00216 (
    .ADR0(id03437),
    .ADR1(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x0 ),
    .ADR2(id03427),
    .O(id03490)
  );

  defparam id00217.INIT = 4'h9;
  LUT2 id00217 (
    .ADR0(id03526),
    .ADR1(id03521),
    .O(id03484)
  );

  defparam id00218.INIT = 16'h9669;
  LUT4 id00218 (
    .ADR0(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x2 ),
    .O(id03526)
  );

  defparam id00219.INIT = 8'hE8;
  LUT3 id00219 (
    .ADR0(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x2 ),
    .O(id03521)
  );

  defparam id00220.INIT = 16'h7117;
  LUT4 id00220 (
    .ADR0(id03433),
    .ADR1(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x0 ),
    .ADR2(id03439),
    .ADR3(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x3 ),
    .O(id03486)
  );

  defparam id00221.INIT = 16'h6996;
  LUT4 id00221 (
    .ADR0(id03514),
    .ADR1(id03528),
    .ADR2(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x3 ),
    .O(id03516)
  );

  defparam id00222.INIT = 4'h6;
  LUT2 id00222 (
    .ADR0(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x2 ),
    .O(id03514)
  );

  defparam id00223.INIT = 8'hE8;
  LUT3 id00223 (
    .ADR0(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x2 ),
    .O(id03528)
  );

  defparam id00224.INIT = 8'hB2;
  LUT3 id00224 (
    .ADR0(id03418),
    .ADR1(id03428),
    .ADR2(id03431),
    .O(id03488)
  );

  defparam id00225.INIT = 8'h35;
  LUT3 id00225 (
    .ADR0(id03480),
    .ADR1(id03445),
    .ADR2(id03435),
    .O(id03545)
  );

  defparam id00226.INIT = 4'h6;
  LUT2 id00226 (
    .ADR0(id03522),
    .ADR1(id03524),
    .O(id03539)
  );

  defparam id00227.INIT = 16'h9669;
  LUT4 id00227 (
    .ADR0(id03534),
    .ADR1(id03536),
    .ADR2(id03530),
    .ADR3(VCC_NET),
    .O(id03522)
  );

  defparam id00228.INIT = 8'h35;
  LUT3 id00228 (
    .ADR0(id03517),
    .ADR1(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x0 ),
    .ADR2(id03482),
    .O(id03534)
  );

  defparam id00229.INIT = 4'h9;
  LUT2 id00229 (
    .ADR0(id03532),
    .ADR1(id03542),
    .O(id03536)
  );

  defparam id00230.INIT = 16'h9669;
  LUT4 id00230 (
    .ADR0(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x2 ),
    .O(id03532)
  );

  defparam id00231.INIT = 8'hE8;
  LUT3 id00231 (
    .ADR0(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x2 ),
    .O(id03542)
  );

  defparam id00232.INIT = 8'h80;
  LUT3 id00232 (
    .ADR0(\u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[38].u_compressor42_cell.x3 ),
    .O(id03530)
  );

  defparam id00233.INIT = 8'hD4;
  LUT3 id00233 (
    .ADR0(id03447),
    .ADR1(id03441),
    .ADR2(id03443),
    .O(id03524)
  );

  defparam id00234.INIT = 4'h1;
  LUT2 id00234 (
    .ADR0(id03529),
    .ADR1(id03523),
    .O(id03187)
  );

  defparam id00235.INIT = 4'h9;
  LUT2 id00235 (
    .ADR0(id03544),
    .ADR1(id03538),
    .O(\net_Buf-pad-result[40] )
  );

  defparam id00236.INIT = 4'h1;
  LUT2 id00236 (
    .ADR0(id03540),
    .ADR1(id03527),
    .O(id03544)
  );

  defparam id00237.INIT = 16'h00D4;
  LUT4 id00237 (
    .ADR0(id03582),
    .ADR1(id03584),
    .ADR2(id03578),
    .ADR3(id03187),
    .O(id03540)
  );

  defparam id00238.INIT = 4'h6;
  LUT2 id00238 (
    .ADR0(id03487),
    .ADR1(id03489),
    .O(id03538)
  );

  defparam id00239.INIT = 4'h4;
  LUT2 id00239 (
    .ADR0(id03525),
    .ADR1(id03535),
    .O(id03487)
  );

  defparam id00240.INIT = 4'h9;
  LUT2 id00240 (
    .ADR0(id03483),
    .ADR1(id03485),
    .O(id03489)
  );

  defparam id00241.INIT = 8'hC5;
  LUT3 id00241 (
    .ADR0(id03539),
    .ADR1(id03537),
    .ADR2(id03531),
    .O(id03483)
  );

  defparam id00242.INIT = 4'h9;
  LUT2 id00242 (
    .ADR0(id03232),
    .ADR1(id03242),
    .O(id03485)
  );

  defparam id00243.INIT = 16'h6996;
  LUT4 id00243 (
    .ADR0(id03236),
    .ADR1(id03231),
    .ADR2(id03244),
    .ADR3(id03238),
    .O(id03232)
  );

  defparam id00244.INIT = 8'hC5;
  LUT3 id00244 (
    .ADR0(id03516),
    .ADR1(id03488),
    .ADR2(id03541),
    .O(id03236)
  );

  defparam id00245.INIT = 4'h9;
  LUT2 id00245 (
    .ADR0(id03243),
    .ADR1(id03245),
    .O(id03231)
  );

  defparam id00246.INIT = 16'h6996;
  LUT4 id00246 (
    .ADR0(id03168),
    .ADR1(id03230),
    .ADR2(id03239),
    .ADR3(id03241),
    .O(id03243)
  );

  defparam id00247.INIT = 8'h35;
  LUT3 id00247 (
    .ADR0(id03521),
    .ADR1(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x0 ),
    .ADR2(id03526),
    .O(id03168)
  );

  defparam id00248.INIT = 4'h9;
  LUT2 id00248 (
    .ADR0(id03186),
    .ADR1(id03247),
    .O(id03230)
  );

  defparam id00249.INIT = 16'h9669;
  LUT4 id00249 (
    .ADR0(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x2 ),
    .O(id03186)
  );

  defparam id00250.INIT = 8'hE8;
  LUT3 id00250 (
    .ADR0(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x2 ),
    .O(id03247)
  );

  defparam id00251.INIT = 16'h7117;
  LUT4 id00251 (
    .ADR0(id03528),
    .ADR1(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x0 ),
    .ADR2(id03514),
    .ADR3(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x3 ),
    .O(id03239)
  );

  defparam id00252.INIT = 16'h6996;
  LUT4 id00252 (
    .ADR0(id03233),
    .ADR1(id03189),
    .ADR2(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x3 ),
    .O(id03241)
  );

  defparam id00253.INIT = 4'h6;
  LUT2 id00253 (
    .ADR0(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x2 ),
    .O(id03233)
  );

  defparam id00254.INIT = 8'hE8;
  LUT3 id00254 (
    .ADR0(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x2 ),
    .O(id03189)
  );

  defparam id00255.INIT = 8'hB2;
  LUT3 id00255 (
    .ADR0(id03490),
    .ADR1(id03484),
    .ADR2(id03486),
    .O(id03245)
  );

  defparam id00256.INIT = 8'h35;
  LUT3 id00256 (
    .ADR0(VCC_NET),
    .ADR1(id03524),
    .ADR2(id03522),
    .O(id03244)
  );

  defparam id00257.INIT = 4'h6;
  LUT2 id00257 (
    .ADR0(id03188),
    .ADR1(id03183),
    .O(id03238)
  );

  defparam id00258.INIT = 16'h53AC;
  LUT4 id00258 (
    .ADR0(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x0 ),
    .ADR1(id03542),
    .ADR2(id03532),
    .ADR3(id03182),
    .O(id03188)
  );

  defparam id00259.INIT = 4'h9;
  LUT2 id00259 (
    .ADR0(id03184),
    .ADR1(id03195),
    .O(id03182)
  );

  defparam id00260.INIT = 16'h9669;
  LUT4 id00260 (
    .ADR0(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x2 ),
    .O(id03184)
  );

  defparam id00261.INIT = 8'hE8;
  LUT3 id00261 (
    .ADR0(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x2 ),
    .O(id03195)
  );

  defparam id00262.INIT = 8'hD4;
  LUT3 id00262 (
    .ADR0(id03534),
    .ADR1(id03536),
    .ADR2(id03530),
    .O(id03183)
  );

  defparam id00263.INIT = 8'hB2;
  LUT3 id00263 (
    .ADR0(id03533),
    .ADR1(id03543),
    .ADR2(id03545),
    .O(id03242)
  );

  defparam id00264.INIT = 16'h2BD4;
  LUT4 id00264 (
    .ADR0(id03544),
    .ADR1(id03487),
    .ADR2(id03489),
    .ADR3(id03194),
    .O(\net_Buf-pad-result[41] )
  );

  defparam id00265.INIT = 4'h6;
  LUT2 id00265 (
    .ADR0(id03197),
    .ADR1(id03196),
    .O(id03194)
  );

  defparam id00266.INIT = 4'h4;
  LUT2 id00266 (
    .ADR0(id03483),
    .ADR1(id03485),
    .O(id03197)
  );

  defparam id00267.INIT = 4'h9;
  LUT2 id00267 (
    .ADR0(id03191),
    .ADR1(id03190),
    .O(id03196)
  );

  defparam id00268.INIT = 8'hC5;
  LUT3 id00268 (
    .ADR0(id03238),
    .ADR1(id03242),
    .ADR2(id03232),
    .O(id03191)
  );

  defparam id00269.INIT = 4'h9;
  LUT2 id00269 (
    .ADR0(id03193),
    .ADR1(id03192),
    .O(id03190)
  );

  defparam id00270.INIT = 16'h9669;
  LUT4 id00270 (
    .ADR0(id03203),
    .ADR1(id03202),
    .ADR2(id03205),
    .ADR3(id03204),
    .O(id03193)
  );

  defparam id00271.INIT = 4'h8;
  LUT2 id00271 (
    .ADR0(id03188),
    .ADR1(id03183),
    .O(id03203)
  );

  defparam id00272.INIT = 8'hC5;
  LUT3 id00272 (
    .ADR0(id03241),
    .ADR1(id03245),
    .ADR2(id03243),
    .O(id03202)
  );

  defparam id00273.INIT = 4'h6;
  LUT2 id00273 (
    .ADR0(id03199),
    .ADR1(id03198),
    .O(id03205)
  );

  defparam id00274.INIT = 16'h9669;
  LUT4 id00274 (
    .ADR0(id03201),
    .ADR1(id03200),
    .ADR2(id03211),
    .ADR3(id03210),
    .O(id03199)
  );

  defparam id00275.INIT = 8'h35;
  LUT3 id00275 (
    .ADR0(id03247),
    .ADR1(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x0 ),
    .ADR2(id03186),
    .O(id03201)
  );

  defparam id00276.INIT = 4'h9;
  LUT2 id00276 (
    .ADR0(id03213),
    .ADR1(id03212),
    .O(id03200)
  );

  defparam id00277.INIT = 16'h9669;
  LUT4 id00277 (
    .ADR0(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x2 ),
    .O(id03213)
  );

  defparam id00278.INIT = 8'hE8;
  LUT3 id00278 (
    .ADR0(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x2 ),
    .O(id03212)
  );

  defparam id00279.INIT = 16'h7117;
  LUT4 id00279 (
    .ADR0(id03189),
    .ADR1(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x0 ),
    .ADR2(id03233),
    .ADR3(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x3 ),
    .O(id03211)
  );

  defparam id00280.INIT = 16'h6996;
  LUT4 id00280 (
    .ADR0(id03207),
    .ADR1(id03206),
    .ADR2(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x3 ),
    .O(id03210)
  );

  defparam id00281.INIT = 4'h6;
  LUT2 id00281 (
    .ADR0(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x2 ),
    .O(id03207)
  );

  defparam id00282.INIT = 8'hE8;
  LUT3 id00282 (
    .ADR0(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x2 ),
    .O(id03206)
  );

  defparam id00283.INIT = 8'hB2;
  LUT3 id00283 (
    .ADR0(id03168),
    .ADR1(id03230),
    .ADR2(id03239),
    .O(id03198)
  );

  defparam id00284.INIT = 4'h6;
  LUT2 id00284 (
    .ADR0(id03209),
    .ADR1(id03208),
    .O(id03204)
  );

  defparam id00285.INIT = 16'hCA00;
  LUT4 id00285 (
    .ADR0(id03542),
    .ADR1(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x0 ),
    .ADR2(id03532),
    .ADR3(id03182),
    .O(id03209)
  );

  defparam id00286.INIT = 16'h53AC;
  LUT4 id00286 (
    .ADR0(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x0 ),
    .ADR1(id03195),
    .ADR2(id03184),
    .ADR3(id03519),
    .O(id03208)
  );

  defparam id00287.INIT = 4'h9;
  LUT2 id00287 (
    .ADR0(id03518),
    .ADR1(id03562),
    .O(id03519)
  );

  defparam id00288.INIT = 16'h9669;
  LUT4 id00288 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x2 ),
    .O(id03518)
  );

  defparam id00289.INIT = 8'hE8;
  LUT3 id00289 (
    .ADR0(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x2 ),
    .O(id03562)
  );

  defparam id00290.INIT = 8'hB2;
  LUT3 id00290 (
    .ADR0(id03236),
    .ADR1(id03231),
    .ADR2(id03244),
    .O(id03192)
  );

  defparam id00291.INIT = 4'h9;
  LUT2 id00291 (
    .ADR0(id03565),
    .ADR1(id03556),
    .O(\net_Buf-pad-result[42] )
  );

  defparam id00292.INIT = 4'h1;
  LUT2 id00292 (
    .ADR0(id03564),
    .ADR1(id03566),
    .O(id03565)
  );

  defparam id00293.INIT = 16'hE000;
  LUT4 id00293 (
    .ADR0(id03527),
    .ADR1(id03540),
    .ADR2(id03538),
    .ADR3(id03194),
    .O(id03564)
  );

  defparam id00294.INIT = 16'hE888;
  LUT4 id00294 (
    .ADR0(id03197),
    .ADR1(id03196),
    .ADR2(id03489),
    .ADR3(id03487),
    .O(id03566)
  );

  defparam id00295.INIT = 4'h6;
  LUT2 id00295 (
    .ADR0(id03569),
    .ADR1(id03568),
    .O(id03556)
  );

  defparam id00296.INIT = 4'h4;
  LUT2 id00296 (
    .ADR0(id03191),
    .ADR1(id03190),
    .O(id03569)
  );

  defparam id00297.INIT = 4'h9;
  LUT2 id00297 (
    .ADR0(id03563),
    .ADR1(id03575),
    .O(id03568)
  );

  defparam id00298.INIT = 8'hC5;
  LUT3 id00298 (
    .ADR0(id03204),
    .ADR1(id03192),
    .ADR2(id03193),
    .O(id03563)
  );

  defparam id00299.INIT = 4'h9;
  LUT2 id00299 (
    .ADR0(id03574),
    .ADR1(id03248),
    .O(id03575)
  );

  defparam id00300.INIT = 16'h6996;
  LUT4 id00300 (
    .ADR0(id03252),
    .ADR1(id03251),
    .ADR2(id03254),
    .ADR3(id03253),
    .O(id03574)
  );

  defparam id00301.INIT = 4'h8;
  LUT2 id00301 (
    .ADR0(id03209),
    .ADR1(id03208),
    .O(id03252)
  );

  defparam id00302.INIT = 8'h3A;
  LUT3 id00302 (
    .ADR0(id03198),
    .ADR1(id03210),
    .ADR2(id03199),
    .O(id03251)
  );

  defparam id00303.INIT = 4'h6;
  LUT2 id00303 (
    .ADR0(id03250),
    .ADR1(id03185),
    .O(id03254)
  );

  defparam id00304.INIT = 16'h9669;
  LUT4 id00304 (
    .ADR0(id03163),
    .ADR1(id03262),
    .ADR2(id03413),
    .ADR3(id03410),
    .O(id03250)
  );

  defparam id00305.INIT = 8'h35;
  LUT3 id00305 (
    .ADR0(id03212),
    .ADR1(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x0 ),
    .ADR2(id03213),
    .O(id03163)
  );

  defparam id00306.INIT = 4'h9;
  LUT2 id00306 (
    .ADR0(id03411),
    .ADR1(id03269),
    .O(id03262)
  );

  defparam id00307.INIT = 16'h9669;
  LUT4 id00307 (
    .ADR0(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x2 ),
    .O(id03411)
  );

  defparam id00308.INIT = 8'hE8;
  LUT3 id00308 (
    .ADR0(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x2 ),
    .O(id03269)
  );

  defparam id00309.INIT = 16'h7117;
  LUT4 id00309 (
    .ADR0(id03206),
    .ADR1(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x0 ),
    .ADR2(id03207),
    .ADR3(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x3 ),
    .O(id03413)
  );

  defparam id00310.INIT = 16'h6996;
  LUT4 id00310 (
    .ADR0(id03271),
    .ADR1(id03265),
    .ADR2(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x3 ),
    .O(id03410)
  );

  defparam id00311.INIT = 4'h6;
  LUT2 id00311 (
    .ADR0(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x2 ),
    .O(id03271)
  );

  defparam id00312.INIT = 8'hE8;
  LUT3 id00312 (
    .ADR0(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x2 ),
    .O(id03265)
  );

  defparam id00313.INIT = 8'hB2;
  LUT3 id00313 (
    .ADR0(id03201),
    .ADR1(id03200),
    .ADR2(id03211),
    .O(id03185)
  );

  defparam id00314.INIT = 4'h6;
  LUT2 id00314 (
    .ADR0(id03412),
    .ADR1(id03277),
    .O(id03253)
  );

  defparam id00315.INIT = 16'hCA00;
  LUT4 id00315 (
    .ADR0(id03195),
    .ADR1(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x0 ),
    .ADR2(id03184),
    .ADR3(id03519),
    .O(id03412)
  );

  defparam id00316.INIT = 16'h53AC;
  LUT4 id00316 (
    .ADR0(VCC_NET),
    .ADR1(id03562),
    .ADR2(id03518),
    .ADR3(id03278),
    .O(id03277)
  );

  defparam id00317.INIT = 16'h17E8;
  LUT4 id00317 (
    .ADR0(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id03273),
    .O(id03278)
  );

  defparam id00318.INIT = 8'h96;
  LUT3 id00318 (
    .ADR0(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x2 ),
    .O(id03273)
  );

  defparam id00319.INIT = 8'hB2;
  LUT3 id00319 (
    .ADR0(id03203),
    .ADR1(id03202),
    .ADR2(id03205),
    .O(id03248)
  );

  defparam id00320.INIT = 16'hD42B;
  LUT4 id00320 (
    .ADR0(id03565),
    .ADR1(id03569),
    .ADR2(id03568),
    .ADR3(id03275),
    .O(\net_Buf-pad-result[43] )
  );

  defparam id00321.INIT = 4'h9;
  LUT2 id00321 (
    .ADR0(id03405),
    .ADR1(id03407),
    .O(id03275)
  );

  defparam id00322.INIT = 4'h4;
  LUT2 id00322 (
    .ADR0(id03563),
    .ADR1(id03575),
    .O(id03405)
  );

  defparam id00323.INIT = 4'h9;
  LUT2 id00323 (
    .ADR0(id03263),
    .ADR1(id03261),
    .O(id03407)
  );

  defparam id00324.INIT = 8'h35;
  LUT3 id00324 (
    .ADR0(id03248),
    .ADR1(id03253),
    .ADR2(id03574),
    .O(id03263)
  );

  defparam id00325.INIT = 4'h9;
  LUT2 id00325 (
    .ADR0(id03409),
    .ADR1(id03270),
    .O(id03261)
  );

  defparam id00326.INIT = 16'h6996;
  LUT4 id00326 (
    .ADR0(id03272),
    .ADR1(id03266),
    .ADR2(id03268),
    .ADR3(id03267),
    .O(id03409)
  );

  defparam id00327.INIT = 4'h8;
  LUT2 id00327 (
    .ADR0(id03412),
    .ADR1(id03277),
    .O(id03272)
  );

  defparam id00328.INIT = 8'h3A;
  LUT3 id00328 (
    .ADR0(id03185),
    .ADR1(id03410),
    .ADR2(id03250),
    .O(id03266)
  );

  defparam id00329.INIT = 4'h9;
  LUT2 id00329 (
    .ADR0(id03279),
    .ADR1(id03274),
    .O(id03268)
  );

  defparam id00330.INIT = 16'h6996;
  LUT4 id00330 (
    .ADR0(id03276),
    .ADR1(id03406),
    .ADR2(id03408),
    .ADR3(id03312),
    .O(id03279)
  );

  defparam id00331.INIT = 8'h35;
  LUT3 id00331 (
    .ADR0(id03269),
    .ADR1(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x0 ),
    .ADR2(id03411),
    .O(id03276)
  );

  defparam id00332.INIT = 4'h9;
  LUT2 id00332 (
    .ADR0(id03476),
    .ADR1(id03477),
    .O(id03406)
  );

  defparam id00333.INIT = 16'h9669;
  LUT4 id00333 (
    .ADR0(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x2 ),
    .O(id03476)
  );

  defparam id00334.INIT = 8'hE8;
  LUT3 id00334 (
    .ADR0(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x2 ),
    .O(id03477)
  );

  defparam id00335.INIT = 16'h7117;
  LUT4 id00335 (
    .ADR0(id03265),
    .ADR1(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x0 ),
    .ADR2(id03271),
    .ADR3(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x3 ),
    .O(id03408)
  );

  defparam id00336.INIT = 16'h6996;
  LUT4 id00336 (
    .ADR0(id03466),
    .ADR1(id03471),
    .ADR2(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x3 ),
    .O(id03312)
  );

  defparam id00337.INIT = 4'h6;
  LUT2 id00337 (
    .ADR0(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x2 ),
    .O(id03466)
  );

  defparam id00338.INIT = 8'hE8;
  LUT3 id00338 (
    .ADR0(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x2 ),
    .O(id03471)
  );

  defparam id00339.INIT = 8'hB2;
  LUT3 id00339 (
    .ADR0(id03163),
    .ADR1(id03262),
    .ADR2(id03413),
    .O(id03274)
  );

  defparam id00340.INIT = 4'h6;
  LUT2 id00340 (
    .ADR0(id03567),
    .ADR1(id03589),
    .O(id03267)
  );

  defparam id00341.INIT = 16'hCA00;
  LUT4 id00341 (
    .ADR0(id03562),
    .ADR1(VCC_NET),
    .ADR2(id03518),
    .ADR3(id03278),
    .O(id03567)
  );

  defparam id00342.INIT = 4'h6;
  LUT2 id00342 (
    .ADR0(id03240),
    .ADR1(id03166),
    .O(id03589)
  );

  defparam id00343.INIT = 16'hE800;
  LUT4 id00343 (
    .ADR0(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id03273),
    .O(id03240)
  );

  defparam id00344.INIT = 16'h6996;
  LUT4 id00344 (
    .ADR0(id03249),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x2 ),
    .O(id03166)
  );

  defparam id00345.INIT = 8'hE8;
  LUT3 id00345 (
    .ADR0(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x2 ),
    .O(id03249)
  );

  defparam id00346.INIT = 8'hB2;
  LUT3 id00346 (
    .ADR0(id03252),
    .ADR1(id03251),
    .ADR2(id03254),
    .O(id03270)
  );

  defparam id00347.INIT = 4'h9;
  LUT2 id00347 (
    .ADR0(id03264),
    .ADR1(id02572),
    .O(\net_Buf-pad-result[44] )
  );

  defparam id00348.INIT = 4'h1;
  LUT2 id00348 (
    .ADR0(id02595),
    .ADR1(id02573),
    .O(id03264)
  );

  defparam id00349.INIT = 16'h0E00;
  LUT4 id00349 (
    .ADR0(id03566),
    .ADR1(id03564),
    .ADR2(id03275),
    .ADR3(id03556),
    .O(id02595)
  );

  defparam id00350.INIT = 16'hB200;
  LUT4 id00350 (
    .ADR0(id03569),
    .ADR1(id03563),
    .ADR2(id03575),
    .ADR3(id03407),
    .O(id02573)
  );

  defparam id00351.INIT = 4'h6;
  LUT2 id00351 (
    .ADR0(id02575),
    .ADR1(id02577),
    .O(id02572)
  );

  defparam id00352.INIT = 4'h4;
  LUT2 id00352 (
    .ADR0(id03263),
    .ADR1(id03261),
    .O(id02575)
  );

  defparam id00353.INIT = 4'h9;
  LUT2 id00353 (
    .ADR0(id02576),
    .ADR1(id02574),
    .O(id02577)
  );

  defparam id00354.INIT = 8'h35;
  LUT3 id00354 (
    .ADR0(id03270),
    .ADR1(id03267),
    .ADR2(id03409),
    .O(id02576)
  );

  defparam id00355.INIT = 4'h6;
  LUT2 id00355 (
    .ADR0(id02827),
    .ADR1(id02829),
    .O(id02574)
  );

  defparam id00356.INIT = 16'h6996;
  LUT4 id00356 (
    .ADR0(id02831),
    .ADR1(id02830),
    .ADR2(id02828),
    .ADR3(id03656),
    .O(id02827)
  );

  defparam id00357.INIT = 4'h8;
  LUT2 id00357 (
    .ADR0(id03567),
    .ADR1(id03589),
    .O(id02831)
  );

  defparam id00358.INIT = 8'hC5;
  LUT3 id00358 (
    .ADR0(id03312),
    .ADR1(id03274),
    .ADR2(id03279),
    .O(id02830)
  );

  defparam id00359.INIT = 4'h9;
  LUT2 id00359 (
    .ADR0(id03637),
    .ADR1(id03639),
    .O(id02828)
  );

  defparam id00360.INIT = 16'h6996;
  LUT4 id00360 (
    .ADR0(id03638),
    .ADR1(id03657),
    .ADR2(id03655),
    .ADR3(id03653),
    .O(id03637)
  );

  defparam id00361.INIT = 8'h35;
  LUT3 id00361 (
    .ADR0(id03477),
    .ADR1(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x0 ),
    .ADR2(id03476),
    .O(id03638)
  );

  defparam id00362.INIT = 4'h9;
  LUT2 id00362 (
    .ADR0(id02819),
    .ADR1(id02818),
    .O(id03657)
  );

  defparam id00363.INIT = 16'h9669;
  LUT4 id00363 (
    .ADR0(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x2 ),
    .O(id02819)
  );

  defparam id00364.INIT = 8'hE8;
  LUT3 id00364 (
    .ADR0(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x2 ),
    .O(id02818)
  );

  defparam id00365.INIT = 16'h7117;
  LUT4 id00365 (
    .ADR0(id03471),
    .ADR1(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x0 ),
    .ADR2(id03466),
    .ADR3(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x3 ),
    .O(id03655)
  );

  defparam id00366.INIT = 16'h6996;
  LUT4 id00366 (
    .ADR0(id02565),
    .ADR1(id02566),
    .ADR2(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x3 ),
    .O(id03653)
  );

  defparam id00367.INIT = 4'h6;
  LUT2 id00367 (
    .ADR0(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x2 ),
    .O(id02565)
  );

  defparam id00368.INIT = 8'hE8;
  LUT3 id00368 (
    .ADR0(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x2 ),
    .O(id02566)
  );

  defparam id00369.INIT = 8'hB2;
  LUT3 id00369 (
    .ADR0(id03276),
    .ADR1(id03406),
    .ADR2(id03408),
    .O(id03639)
  );

  defparam id00370.INIT = 8'hE1;
  LUT3 id00370 (
    .ADR0(id02571),
    .ADR1(id02568),
    .ADR2(id02567),
    .O(id03656)
  );

  defparam id00371.INIT = 4'h8;
  LUT2 id00371 (
    .ADR0(id03240),
    .ADR1(id03166),
    .O(id02571)
  );

  defparam id00372.INIT = 16'h9600;
  LUT4 id00372 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x2 ),
    .ADR3(id03249),
    .O(id02568)
  );

  defparam id00373.INIT = 8'h96;
  LUT3 id00373 (
    .ADR0(id02570),
    .ADR1(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 ),
    .O(id02567)
  );

  defparam id00374.INIT = 8'hE8;
  LUT3 id00374 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x2 ),
    .O(id02570)
  );

  defparam id00375.INIT = 8'hB2;
  LUT3 id00375 (
    .ADR0(id03272),
    .ADR1(id03266),
    .ADR2(id03268),
    .O(id02829)
  );

  defparam id00376.INIT = 16'h2BD4;
  LUT4 id00376 (
    .ADR0(id03264),
    .ADR1(id02575),
    .ADR2(id02577),
    .ADR3(id02569),
    .O(\net_Buf-pad-result[45] )
  );

  defparam id00377.INIT = 4'h6;
  LUT2 id00377 (
    .ADR0(id02826),
    .ADR1(id02823),
    .O(id02569)
  );

  defparam id00378.INIT = 4'h4;
  LUT2 id00378 (
    .ADR0(id02576),
    .ADR1(id02574),
    .O(id02826)
  );

  defparam id00379.INIT = 4'h9;
  LUT2 id00379 (
    .ADR0(id02822),
    .ADR1(id02825),
    .O(id02823)
  );

  defparam id00380.INIT = 8'h3A;
  LUT3 id00380 (
    .ADR0(id03656),
    .ADR1(id02829),
    .ADR2(id02827),
    .O(id02822)
  );

  defparam id00381.INIT = 4'h6;
  LUT2 id00381 (
    .ADR0(id02824),
    .ADR1(id03633),
    .O(id02825)
  );

  defparam id00382.INIT = 16'h6996;
  LUT4 id00382 (
    .ADR0(id03635),
    .ADR1(id03634),
    .ADR2(id03632),
    .ADR3(id03636),
    .O(id02824)
  );

  defparam id00383.INIT = 8'hC5;
  LUT3 id00383 (
    .ADR0(id03653),
    .ADR1(id03639),
    .ADR2(id03637),
    .O(id03635)
  );

  defparam id00384.INIT = 4'h6;
  LUT2 id00384 (
    .ADR0(id03641),
    .ADR1(id03642),
    .O(id03634)
  );

  defparam id00385.INIT = 16'h9669;
  LUT4 id00385 (
    .ADR0(id02820),
    .ADR1(id02821),
    .ADR2(id02584),
    .ADR3(id02583),
    .O(id03641)
  );

  defparam id00386.INIT = 8'h35;
  LUT3 id00386 (
    .ADR0(id02818),
    .ADR1(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x0 ),
    .ADR2(id02819),
    .O(id02820)
  );

  defparam id00387.INIT = 4'h9;
  LUT2 id00387 (
    .ADR0(id02578),
    .ADR1(id02580),
    .O(id02821)
  );

  defparam id00388.INIT = 16'h9669;
  LUT4 id00388 (
    .ADR0(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x2 ),
    .O(id02578)
  );

  defparam id00389.INIT = 8'hE8;
  LUT3 id00389 (
    .ADR0(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x2 ),
    .O(id02580)
  );

  defparam id00390.INIT = 16'h7117;
  LUT4 id00390 (
    .ADR0(id02566),
    .ADR1(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x0 ),
    .ADR2(id02565),
    .ADR3(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x3 ),
    .O(id02584)
  );

  defparam id00391.INIT = 16'h6996;
  LUT4 id00391 (
    .ADR0(id02582),
    .ADR1(id02581),
    .ADR2(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x3 ),
    .O(id02583)
  );

  defparam id00392.INIT = 4'h6;
  LUT2 id00392 (
    .ADR0(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x2 ),
    .O(id02582)
  );

  defparam id00393.INIT = 8'hE8;
  LUT3 id00393 (
    .ADR0(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x2 ),
    .O(id02581)
  );

  defparam id00394.INIT = 8'hB2;
  LUT3 id00394 (
    .ADR0(id03638),
    .ADR1(id03657),
    .ADR2(id03655),
    .O(id03642)
  );

  defparam id00395.INIT = 4'h8;
  LUT2 id00395 (
    .ADR0(id02571),
    .ADR1(id02567),
    .O(id03632)
  );

  defparam id00396.INIT = 16'hF807;
  LUT4 id00396 (
    .ADR0(id02568),
    .ADR1(id02567),
    .ADR2(id02579),
    .ADR3(id02804),
    .O(id03636)
  );

  defparam id00397.INIT = 8'h60;
  LUT3 id00397 (
    .ADR0(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(id02570),
    .O(id02579)
  );

  defparam id00398.INIT = 16'h8778;
  LUT4 id00398 (
    .ADR0(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(\u_compressor42_l0_1.CELLS[39].u_compressor42_cell.x3 ),
    .ADR3(VCC_NET),
    .O(id02804)
  );

  defparam id00399.INIT = 8'hB2;
  LUT3 id00399 (
    .ADR0(id02831),
    .ADR1(id02830),
    .ADR2(id02828),
    .O(id03633)
  );

  defparam id00400.INIT = 4'h9;
  LUT2 id00400 (
    .ADR0(id02797),
    .ADR1(id02799),
    .O(\net_Buf-pad-result[46] )
  );

  defparam id00401.INIT = 4'h4;
  LUT2 id00401 (
    .ADR0(id02798),
    .ADR1(id02805),
    .O(id02797)
  );

  defparam id00402.INIT = 16'hE000;
  LUT4 id00402 (
    .ADR0(id02573),
    .ADR1(id02595),
    .ADR2(id02572),
    .ADR3(id02569),
    .O(id02798)
  );

  defparam id00403.INIT = 16'h07FF;
  LUT4 id00403 (
    .ADR0(id02575),
    .ADR1(id02577),
    .ADR2(id02826),
    .ADR3(id02823),
    .O(id02805)
  );

  defparam id00404.INIT = 4'h6;
  LUT2 id00404 (
    .ADR0(id03650),
    .ADR1(id03649),
    .O(id02799)
  );

  defparam id00405.INIT = 4'h4;
  LUT2 id00405 (
    .ADR0(id02822),
    .ADR1(id02825),
    .O(id03650)
  );

  defparam id00406.INIT = 4'h6;
  LUT2 id00406 (
    .ADR0(id03652),
    .ADR1(id03651),
    .O(id03649)
  );

  defparam id00407.INIT = 4'h6;
  LUT2 id00407 (
    .ADR0(id03645),
    .ADR1(id03647),
    .O(id03652)
  );

  defparam id00408.INIT = 16'h6996;
  LUT4 id00408 (
    .ADR0(id02803),
    .ADR1(id02802),
    .ADR2(id02546),
    .ADR3(id02547),
    .O(id03645)
  );

  defparam id00409.INIT = 8'h3A;
  LUT3 id00409 (
    .ADR0(id03642),
    .ADR1(id02583),
    .ADR2(id03641),
    .O(id02803)
  );

  defparam id00410.INIT = 4'h9;
  LUT2 id00410 (
    .ADR0(id02549),
    .ADR1(id02551),
    .O(id02802)
  );

  defparam id00411.INIT = 16'h6996;
  LUT4 id00411 (
    .ADR0(id02550),
    .ADR1(id02548),
    .ADR2(id02552),
    .ADR3(id02814),
    .O(id02549)
  );

  defparam id00412.INIT = 8'h35;
  LUT3 id00412 (
    .ADR0(id02580),
    .ADR1(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x0 ),
    .ADR2(id02578),
    .O(id02550)
  );

  defparam id00413.INIT = 4'h9;
  LUT2 id00413 (
    .ADR0(id02816),
    .ADR1(id02815),
    .O(id02548)
  );

  defparam id00414.INIT = 16'h9669;
  LUT4 id00414 (
    .ADR0(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x2 ),
    .O(id02816)
  );

  defparam id00415.INIT = 8'hE8;
  LUT3 id00415 (
    .ADR0(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x2 ),
    .O(id02815)
  );

  defparam id00416.INIT = 16'h7117;
  LUT4 id00416 (
    .ADR0(id02581),
    .ADR1(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x0 ),
    .ADR2(id02582),
    .ADR3(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x3 ),
    .O(id02552)
  );

  defparam id00417.INIT = 16'h6996;
  LUT4 id00417 (
    .ADR0(id02813),
    .ADR1(id02817),
    .ADR2(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x3 ),
    .O(id02814)
  );

  defparam id00418.INIT = 4'h6;
  LUT2 id00418 (
    .ADR0(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x2 ),
    .O(id02813)
  );

  defparam id00419.INIT = 8'hE8;
  LUT3 id00419 (
    .ADR0(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x2 ),
    .O(id02817)
  );

  defparam id00420.INIT = 8'hB2;
  LUT3 id00420 (
    .ADR0(id02820),
    .ADR1(id02821),
    .ADR2(id02584),
    .O(id02551)
  );

  defparam id00421.INIT = 8'h80;
  LUT3 id00421 (
    .ADR0(id02568),
    .ADR1(id02567),
    .ADR2(id02804),
    .O(id02546)
  );

  defparam id00422.INIT = 16'h7887;
  LUT4 id00422 (
    .ADR0(id02579),
    .ADR1(id02804),
    .ADR2(id03623),
    .ADR3(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ),
    .O(id02547)
  );

  defparam id00423.INIT = 4'h1;
  LUT2 id00423 (
    .ADR0(id03624),
    .ADR1(id03622),
    .O(id03623)
  );

  defparam id00424.INIT = 4'h8;
  LUT2 id00424 (
    .ADR0(\u_compressor42_l0_1.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .O(id03624)
  );

  defparam id00425.INIT = 16'h6000;
  LUT4 id00425 (
    .ADR0(\u_compressor42_l0_1.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 ),
    .O(id03622)
  );

  defparam id00426.INIT = 8'hD4;
  LUT3 id00426 (
    .ADR0(id03635),
    .ADR1(id03634),
    .ADR2(id03632),
    .O(id03647)
  );

  defparam id00427.INIT = 8'h3A;
  LUT3 id00427 (
    .ADR0(id03636),
    .ADR1(id03633),
    .ADR2(id02824),
    .O(id03651)
  );

  defparam id00428.INIT = 16'hD42B;
  LUT4 id00428 (
    .ADR0(id02797),
    .ADR1(id03650),
    .ADR2(id03649),
    .ADR3(id03621),
    .O(\net_Buf-pad-result[47] )
  );

  defparam id00429.INIT = 4'h9;
  LUT2 id00429 (
    .ADR0(id02800),
    .ADR1(id02801),
    .O(id03621)
  );

  defparam id00430.INIT = 4'h1;
  LUT2 id00430 (
    .ADR0(id03652),
    .ADR1(id03651),
    .O(id02800)
  );

  defparam id00431.INIT = 4'h6;
  LUT2 id00431 (
    .ADR0(id02544),
    .ADR1(id02545),
    .O(id02801)
  );

  defparam id00432.INIT = 4'h9;
  LUT2 id00432 (
    .ADR0(id02561),
    .ADR1(id02563),
    .O(id02544)
  );

  defparam id00433.INIT = 16'h6996;
  LUT4 id00433 (
    .ADR0(id02560),
    .ADR1(id02564),
    .ADR2(id02562),
    .ADR3(id02809),
    .O(id02561)
  );

  defparam id00434.INIT = 8'hC5;
  LUT3 id00434 (
    .ADR0(id02814),
    .ADR1(id02551),
    .ADR2(id02549),
    .O(id02560)
  );

  defparam id00435.INIT = 4'h6;
  LUT2 id00435 (
    .ADR0(id02811),
    .ADR1(id02808),
    .O(id02564)
  );

  defparam id00436.INIT = 16'h9669;
  LUT4 id00436 (
    .ADR0(id02812),
    .ADR1(id02810),
    .ADR2(id02806),
    .ADR3(id02807),
    .O(id02811)
  );

  defparam id00437.INIT = 8'h35;
  LUT3 id00437 (
    .ADR0(id02815),
    .ADR1(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x0 ),
    .ADR2(id02816),
    .O(id02812)
  );

  defparam id00438.INIT = 4'h9;
  LUT2 id00438 (
    .ADR0(id02553),
    .ADR1(id02554),
    .O(id02810)
  );

  defparam id00439.INIT = 16'h9669;
  LUT4 id00439 (
    .ADR0(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x2 ),
    .O(id02553)
  );

  defparam id00440.INIT = 8'hE8;
  LUT3 id00440 (
    .ADR0(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x2 ),
    .O(id02554)
  );

  defparam id00441.INIT = 16'h7117;
  LUT4 id00441 (
    .ADR0(id02817),
    .ADR1(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x0 ),
    .ADR2(id02813),
    .ADR3(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x3 ),
    .O(id02806)
  );

  defparam id00442.INIT = 16'h6996;
  LUT4 id00442 (
    .ADR0(id02557),
    .ADR1(id02559),
    .ADR2(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x3 ),
    .O(id02807)
  );

  defparam id00443.INIT = 4'h6;
  LUT2 id00443 (
    .ADR0(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x2 ),
    .O(id02557)
  );

  defparam id00444.INIT = 8'hE8;
  LUT3 id00444 (
    .ADR0(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x2 ),
    .O(id02559)
  );

  defparam id00445.INIT = 8'hB2;
  LUT3 id00445 (
    .ADR0(id02550),
    .ADR1(id02548),
    .ADR2(id02552),
    .O(id02808)
  );

  defparam id00446.INIT = 8'h80;
  LUT3 id00446 (
    .ADR0(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ),
    .ADR1(id02804),
    .ADR2(id02579),
    .O(id02562)
  );

  defparam id00447.INIT = 16'hD728;
  LUT4 id00447 (
    .ADR0(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ),
    .ADR1(id03624),
    .ADR2(id03622),
    .ADR3(VCC_NET),
    .O(id02809)
  );

  defparam id00448.INIT = 8'hD4;
  LUT3 id00448 (
    .ADR0(id02803),
    .ADR1(id02802),
    .ADR2(id02546),
    .O(id02563)
  );

  defparam id00449.INIT = 8'hCA;
  LUT3 id00449 (
    .ADR0(id03647),
    .ADR1(id02547),
    .ADR2(id03645),
    .O(id02545)
  );

  defparam id00450.INIT = 16'hE11E;
  LUT4 id00450 (
    .ADR0(id02558),
    .ADR1(id02556),
    .ADR2(id02555),
    .ADR3(id02786),
    .O(\net_Buf-pad-result[48] )
  );

  defparam id00451.INIT = 16'h0D00;
  LUT4 id00451 (
    .ADR0(id02805),
    .ADR1(id02798),
    .ADR2(id03621),
    .ADR3(id02799),
    .O(id02558)
  );

  defparam id00452.INIT = 16'h2B00;
  LUT4 id00452 (
    .ADR0(id03650),
    .ADR1(id03652),
    .ADR2(id03651),
    .ADR3(id02801),
    .O(id02556)
  );

  defparam id00453.INIT = 4'h8;
  LUT2 id00453 (
    .ADR0(id02544),
    .ADR1(id02545),
    .O(id02555)
  );

  defparam id00454.INIT = 4'h9;
  LUT2 id00454 (
    .ADR0(id02788),
    .ADR1(id02787),
    .O(id02786)
  );

  defparam id00455.INIT = 8'h35;
  LUT3 id00455 (
    .ADR0(id02563),
    .ADR1(id02809),
    .ADR2(id02561),
    .O(id02788)
  );

  defparam id00456.INIT = 16'hE11E;
  LUT4 id00456 (
    .ADR0(id02785),
    .ADR1(id02784),
    .ADR2(id03181),
    .ADR3(id03179),
    .O(id02787)
  );

  defparam id00457.INIT = 8'hD4;
  LUT3 id00457 (
    .ADR0(id02560),
    .ADR1(id02564),
    .ADR2(id02562),
    .O(id03181)
  );

  defparam id00458.INIT = 4'h9;
  LUT2 id00458 (
    .ADR0(id03154),
    .ADR1(id03161),
    .O(id03179)
  );

  defparam id00459.INIT = 8'h3A;
  LUT3 id00459 (
    .ADR0(id02808),
    .ADR1(id02807),
    .ADR2(id02811),
    .O(id03154)
  );

  defparam id00460.INIT = 4'h9;
  LUT2 id00460 (
    .ADR0(id02789),
    .ADR1(id02790),
    .O(id03161)
  );

  defparam id00461.INIT = 16'h6996;
  LUT4 id00461 (
    .ADR0(id02526),
    .ADR1(id02525),
    .ADR2(id02530),
    .ADR3(id02527),
    .O(id02789)
  );

  defparam id00462.INIT = 8'h35;
  LUT3 id00462 (
    .ADR0(id02554),
    .ADR1(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x0 ),
    .ADR2(id02553),
    .O(id02526)
  );

  defparam id00463.INIT = 4'h9;
  LUT2 id00463 (
    .ADR0(id02529),
    .ADR1(id02528),
    .O(id02525)
  );

  defparam id00464.INIT = 16'h9669;
  LUT4 id00464 (
    .ADR0(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x2 ),
    .O(id02529)
  );

  defparam id00465.INIT = 8'hE8;
  LUT3 id00465 (
    .ADR0(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x2 ),
    .O(id02528)
  );

  defparam id00466.INIT = 16'h7117;
  LUT4 id00466 (
    .ADR0(id02559),
    .ADR1(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x0 ),
    .ADR2(id02557),
    .ADR3(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x3 ),
    .O(id02530)
  );

  defparam id00467.INIT = 16'h6996;
  LUT4 id00467 (
    .ADR0(id02531),
    .ADR1(id02795),
    .ADR2(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x3 ),
    .O(id02527)
  );

  defparam id00468.INIT = 4'h6;
  LUT2 id00468 (
    .ADR0(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x2 ),
    .O(id02531)
  );

  defparam id00469.INIT = 8'hE8;
  LUT3 id00469 (
    .ADR0(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x2 ),
    .O(id02795)
  );

  defparam id00470.INIT = 8'hB2;
  LUT3 id00470 (
    .ADR0(id02812),
    .ADR1(id02810),
    .ADR2(id02806),
    .O(id02790)
  );

  defparam id00471.INIT = 8'h80;
  LUT3 id00471 (
    .ADR0(id03624),
    .ADR1(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ),
    .ADR2(VCC_NET),
    .O(id02785)
  );

  defparam id00472.INIT = 8'h80;
  LUT3 id00472 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 ),
    .ADR2(id03622),
    .O(id02784)
  );

  defparam id00473.INIT = 8'h69;
  LUT3 id00473 (
    .ADR0(id02794),
    .ADR1(id02793),
    .ADR2(id02796),
    .O(\net_Buf-pad-result[49] )
  );

  defparam id00474.INIT = 16'h1117;
  LUT4 id00474 (
    .ADR0(id02555),
    .ADR1(id02786),
    .ADR2(id02558),
    .ADR3(id02556),
    .O(id02794)
  );

  defparam id00475.INIT = 4'h4;
  LUT2 id00475 (
    .ADR0(id02788),
    .ADR1(id02787),
    .O(id02793)
  );

  defparam id00476.INIT = 4'h9;
  LUT2 id00476 (
    .ADR0(id02979),
    .ADR1(id02978),
    .O(id02796)
  );

  defparam id00477.INIT = 16'h0D57;
  LUT4 id00477 (
    .ADR0(id03181),
    .ADR1(id02784),
    .ADR2(id02785),
    .ADR3(id03179),
    .O(id02979)
  );

  defparam id00478.INIT = 4'h6;
  LUT2 id00478 (
    .ADR0(id02792),
    .ADR1(id02791),
    .O(id02978)
  );

  defparam id00479.INIT = 4'h9;
  LUT2 id00479 (
    .ADR0(id02523),
    .ADR1(id02524),
    .O(id02792)
  );

  defparam id00480.INIT = 8'hC5;
  LUT3 id00480 (
    .ADR0(id02527),
    .ADR1(id02790),
    .ADR2(id02789),
    .O(id02523)
  );

  defparam id00481.INIT = 4'h6;
  LUT2 id00481 (
    .ADR0(id02541),
    .ADR1(id02543),
    .O(id02524)
  );

  defparam id00482.INIT = 16'h9669;
  LUT4 id00482 (
    .ADR0(id02542),
    .ADR1(id02540),
    .ADR2(id02539),
    .ADR3(id02533),
    .O(id02541)
  );

  defparam id00483.INIT = 8'h35;
  LUT3 id00483 (
    .ADR0(id02528),
    .ADR1(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x0 ),
    .ADR2(id02529),
    .O(id02542)
  );

  defparam id00484.INIT = 4'h9;
  LUT2 id00484 (
    .ADR0(id02532),
    .ADR1(id02534),
    .O(id02540)
  );

  defparam id00485.INIT = 16'h9669;
  LUT4 id00485 (
    .ADR0(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x2 ),
    .O(id02532)
  );

  defparam id00486.INIT = 8'hE8;
  LUT3 id00486 (
    .ADR0(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x2 ),
    .O(id02534)
  );

  defparam id00487.INIT = 16'h7117;
  LUT4 id00487 (
    .ADR0(id02795),
    .ADR1(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x0 ),
    .ADR2(id02531),
    .ADR3(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x3 ),
    .O(id02539)
  );

  defparam id00488.INIT = 16'h6996;
  LUT4 id00488 (
    .ADR0(id02536),
    .ADR1(id02538),
    .ADR2(VCC_NET),
    .ADR3(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 ),
    .O(id02533)
  );

  defparam id00489.INIT = 4'h6;
  LUT2 id00489 (
    .ADR0(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x2 ),
    .O(id02536)
  );

  defparam id00490.INIT = 8'hE8;
  LUT3 id00490 (
    .ADR0(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x2 ),
    .O(id02538)
  );

  defparam id00491.INIT = 8'hB2;
  LUT3 id00491 (
    .ADR0(id02526),
    .ADR1(id02525),
    .ADR2(id02530),
    .O(id02543)
  );

  defparam id00492.INIT = 8'hD4;
  LUT3 id00492 (
    .ADR0(id03154),
    .ADR1(id03161),
    .ADR2(id02784),
    .O(id02791)
  );

  defparam id00493.INIT = 16'h2BD4;
  LUT4 id00493 (
    .ADR0(id02794),
    .ADR1(id02793),
    .ADR2(id02796),
    .ADR3(id02537),
    .O(\net_Buf-pad-result[50] )
  );

  defparam id00494.INIT = 4'h6;
  LUT2 id00494 (
    .ADR0(id02535),
    .ADR1(id02497),
    .O(id02537)
  );

  defparam id00495.INIT = 4'h4;
  LUT2 id00495 (
    .ADR0(id02979),
    .ADR1(id02978),
    .O(id02535)
  );

  defparam id00496.INIT = 4'h6;
  LUT2 id00496 (
    .ADR0(id02498),
    .ADR1(id02496),
    .O(id02497)
  );

  defparam id00497.INIT = 4'h8;
  LUT2 id00497 (
    .ADR0(id02792),
    .ADR1(id02791),
    .O(id02498)
  );

  defparam id00498.INIT = 4'h6;
  LUT2 id00498 (
    .ADR0(id02493),
    .ADR1(id02492),
    .O(id02496)
  );

  defparam id00499.INIT = 4'h4;
  LUT2 id00499 (
    .ADR0(id02523),
    .ADR1(id02524),
    .O(id02493)
  );

  defparam id00500.INIT = 4'h9;
  LUT2 id00500 (
    .ADR0(id02495),
    .ADR1(id02494),
    .O(id02492)
  );

  defparam id00501.INIT = 8'h3A;
  LUT3 id00501 (
    .ADR0(id02543),
    .ADR1(id02533),
    .ADR2(id02541),
    .O(id02495)
  );

  defparam id00502.INIT = 4'h9;
  LUT2 id00502 (
    .ADR0(id02507),
    .ADR1(id02506),
    .O(id02494)
  );

  defparam id00503.INIT = 16'h9669;
  LUT4 id00503 (
    .ADR0(id02508),
    .ADR1(id02510),
    .ADR2(id02512),
    .ADR3(id02511),
    .O(id02507)
  );

  defparam id00504.INIT = 8'h35;
  LUT3 id00504 (
    .ADR0(id02534),
    .ADR1(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x0 ),
    .ADR2(id02532),
    .O(id02508)
  );

  defparam id00505.INIT = 4'h9;
  LUT2 id00505 (
    .ADR0(id02509),
    .ADR1(id02499),
    .O(id02510)
  );

  defparam id00506.INIT = 16'h9669;
  LUT4 id00506 (
    .ADR0(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x2 ),
    .O(id02509)
  );

  defparam id00507.INIT = 8'hE8;
  LUT3 id00507 (
    .ADR0(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x2 ),
    .O(id02499)
  );

  defparam id00508.INIT = 16'h7117;
  LUT4 id00508 (
    .ADR0(id02538),
    .ADR1(VCC_NET),
    .ADR2(id02536),
    .ADR3(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 ),
    .O(id02512)
  );

  defparam id00509.INIT = 16'h17E8;
  LUT4 id00509 (
    .ADR0(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id02500),
    .O(id02511)
  );

  defparam id00510.INIT = 8'h96;
  LUT3 id00510 (
    .ADR0(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x2 ),
    .O(id02500)
  );

  defparam id00511.INIT = 8'h71;
  LUT3 id00511 (
    .ADR0(id02542),
    .ADR1(id02539),
    .ADR2(id02540),
    .O(id02506)
  );

  defparam id00512.INIT = 8'h1E;
  LUT3 id00512 (
    .ADR0(id02502),
    .ADR1(id02504),
    .ADR2(id02503),
    .O(\net_Buf-pad-result[51] )
  );

  defparam id00513.INIT = 16'hD400;
  LUT4 id00513 (
    .ADR0(id02794),
    .ADR1(id02793),
    .ADR2(id02796),
    .ADR3(id02537),
    .O(id02502)
  );

  defparam id00514.INIT = 4'h1;
  LUT2 id00514 (
    .ADR0(id02501),
    .ADR1(id02505),
    .O(id02503)
  );

  defparam id00515.INIT = 4'h8;
  LUT2 id00515 (
    .ADR0(id02481),
    .ADR1(id02482),
    .O(id02501)
  );

  defparam id00516.INIT = 4'h8;
  LUT2 id00516 (
    .ADR0(id02498),
    .ADR1(id02496),
    .O(id02481)
  );

  defparam id00517.INIT = 4'h6;
  LUT2 id00517 (
    .ADR0(id02477),
    .ADR1(id02479),
    .O(id02482)
  );

  defparam id00518.INIT = 4'h4;
  LUT2 id00518 (
    .ADR0(id02495),
    .ADR1(id02494),
    .O(id02477)
  );

  defparam id00519.INIT = 4'h9;
  LUT2 id00519 (
    .ADR0(id02476),
    .ADR1(id02480),
    .O(id02479)
  );

  defparam id00520.INIT = 8'h35;
  LUT3 id00520 (
    .ADR0(id02506),
    .ADR1(id02511),
    .ADR2(id02507),
    .O(id02476)
  );

  defparam id00521.INIT = 4'h6;
  LUT2 id00521 (
    .ADR0(id02478),
    .ADR1(id02485),
    .O(id02480)
  );

  defparam id00522.INIT = 16'h6996;
  LUT4 id00522 (
    .ADR0(id02486),
    .ADR1(id02489),
    .ADR2(id02491),
    .ADR3(id02490),
    .O(id02478)
  );

  defparam id00523.INIT = 16'hE800;
  LUT4 id00523 (
    .ADR0(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id02500),
    .O(id02486)
  );

  defparam id00524.INIT = 8'h35;
  LUT3 id00524 (
    .ADR0(id02499),
    .ADR1(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x0 ),
    .ADR2(id02509),
    .O(id02489)
  );

  defparam id00525.INIT = 4'h9;
  LUT2 id00525 (
    .ADR0(id02488),
    .ADR1(id02487),
    .O(id02491)
  );

  defparam id00526.INIT = 16'h9669;
  LUT4 id00526 (
    .ADR0(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x2 ),
    .O(id02488)
  );

  defparam id00527.INIT = 8'hE8;
  LUT3 id00527 (
    .ADR0(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x2 ),
    .O(id02487)
  );

  defparam id00528.INIT = 16'h6996;
  LUT4 id00528 (
    .ADR0(id03178),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x2 ),
    .O(id02490)
  );

  defparam id00529.INIT = 8'hE8;
  LUT3 id00529 (
    .ADR0(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x2 ),
    .O(id03178)
  );

  defparam id00530.INIT = 8'hB2;
  LUT3 id00530 (
    .ADR0(id02508),
    .ADR1(id02510),
    .ADR2(id02512),
    .O(id02485)
  );

  defparam id00531.INIT = 8'h41;
  LUT3 id00531 (
    .ADR0(id02481),
    .ADR1(id03156),
    .ADR2(id02482),
    .O(id02505)
  );

  defparam id00532.INIT = 4'h8;
  LUT2 id00532 (
    .ADR0(id02493),
    .ADR1(id02492),
    .O(id03156)
  );

  defparam id00533.INIT = 4'h8;
  LUT2 id00533 (
    .ADR0(id02535),
    .ADR1(id02497),
    .O(id02504)
  );

  defparam id00534.INIT = 16'h708F;
  LUT4 id00534 (
    .ADR0(id02502),
    .ADR1(id02503),
    .ADR2(id03155),
    .ADR3(id03158),
    .O(\net_Buf-pad-result[52] )
  );

  defparam id00535.INIT = 8'h0B;
  LUT3 id00535 (
    .ADR0(id02505),
    .ADR1(id02504),
    .ADR2(id02501),
    .O(id03155)
  );

  defparam id00536.INIT = 4'h6;
  LUT2 id00536 (
    .ADR0(id02484),
    .ADR1(id02483),
    .O(id03158)
  );

  defparam id00537.INIT = 4'h8;
  LUT2 id00537 (
    .ADR0(id03156),
    .ADR1(id02482),
    .O(id02484)
  );

  defparam id00538.INIT = 4'h6;
  LUT2 id00538 (
    .ADR0(id02474),
    .ADR1(id02473),
    .O(id02483)
  );

  defparam id00539.INIT = 4'h8;
  LUT2 id00539 (
    .ADR0(id02477),
    .ADR1(id02479),
    .O(id02474)
  );

  defparam id00540.INIT = 4'h6;
  LUT2 id00540 (
    .ADR0(id02472),
    .ADR1(id02475),
    .O(id02473)
  );

  defparam id00541.INIT = 4'h4;
  LUT2 id00541 (
    .ADR0(id02476),
    .ADR1(id02480),
    .O(id02472)
  );

  defparam id00542.INIT = 4'h9;
  LUT2 id00542 (
    .ADR0(id02429),
    .ADR1(id02428),
    .O(id02475)
  );

  defparam id00543.INIT = 8'h3A;
  LUT3 id00543 (
    .ADR0(id02485),
    .ADR1(id02490),
    .ADR2(id02478),
    .O(id02429)
  );

  defparam id00544.INIT = 4'h9;
  LUT2 id00544 (
    .ADR0(id02430),
    .ADR1(id02432),
    .O(id02428)
  );

  defparam id00545.INIT = 16'h6996;
  LUT4 id00545 (
    .ADR0(id02434),
    .ADR1(id02433),
    .ADR2(id02431),
    .ADR3(id03085),
    .O(id02430)
  );

  defparam id00546.INIT = 16'h9600;
  LUT4 id00546 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x2 ),
    .ADR3(id03178),
    .O(id02434)
  );

  defparam id00547.INIT = 8'h35;
  LUT3 id00547 (
    .ADR0(id02487),
    .ADR1(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x0 ),
    .ADR2(id02488),
    .O(id02433)
  );

  defparam id00548.INIT = 4'h9;
  LUT2 id00548 (
    .ADR0(id03086),
    .ADR1(id02421),
    .O(id02431)
  );

  defparam id00549.INIT = 16'h9669;
  LUT4 id00549 (
    .ADR0(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x2 ),
    .O(id03086)
  );

  defparam id00550.INIT = 8'hE8;
  LUT3 id00550 (
    .ADR0(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x2 ),
    .O(id02421)
  );

  defparam id00551.INIT = 8'h96;
  LUT3 id00551 (
    .ADR0(id02422),
    .ADR1(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 ),
    .O(id03085)
  );

  defparam id00552.INIT = 8'hE8;
  LUT3 id00552 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x2 ),
    .O(id02422)
  );

  defparam id00553.INIT = 8'hB2;
  LUT3 id00553 (
    .ADR0(id02486),
    .ADR1(id02489),
    .ADR2(id02491),
    .O(id02432)
  );

  defparam id00554.INIT = 8'h1E;
  LUT3 id00554 (
    .ADR0(id02424),
    .ADR1(id02426),
    .ADR2(id02425),
    .O(\net_Buf-pad-result[53] )
  );

  defparam id00555.INIT = 16'h8F00;
  LUT4 id00555 (
    .ADR0(id02503),
    .ADR1(id02502),
    .ADR2(id03155),
    .ADR3(id03158),
    .O(id02424)
  );

  defparam id00556.INIT = 4'h6;
  LUT2 id00556 (
    .ADR0(id02423),
    .ADR1(id02427),
    .O(id02425)
  );

  defparam id00557.INIT = 4'h6;
  LUT2 id00557 (
    .ADR0(id02440),
    .ADR1(id02441),
    .O(id02423)
  );

  defparam id00558.INIT = 4'h6;
  LUT2 id00558 (
    .ADR0(id02436),
    .ADR1(id02438),
    .O(id02440)
  );

  defparam id00559.INIT = 4'h9;
  LUT2 id00559 (
    .ADR0(id02435),
    .ADR1(id02439),
    .O(id02436)
  );

  defparam id00560.INIT = 4'h6;
  LUT2 id00560 (
    .ADR0(id02437),
    .ADR1(id02402),
    .O(id02435)
  );

  defparam id00561.INIT = 8'h69;
  LUT3 id00561 (
    .ADR0(id02403),
    .ADR1(id02406),
    .ADR2(id02408),
    .O(id02437)
  );

  defparam id00562.INIT = 4'h6;
  LUT2 id00562 (
    .ADR0(id02407),
    .ADR1(id02405),
    .O(id02403)
  );

  defparam id00563.INIT = 8'h60;
  LUT3 id00563 (
    .ADR0(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(id02422),
    .O(id02405)
  );

  defparam id00564.INIT = 16'h8778;
  LUT4 id00564 (
    .ADR0(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(\u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 ),
    .ADR3(VCC_NET),
    .O(id02407)
  );

  defparam id00565.INIT = 8'h35;
  LUT3 id00565 (
    .ADR0(id02421),
    .ADR1(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x0 ),
    .ADR2(id03086),
    .O(id02406)
  );

  defparam id00566.INIT = 4'h9;
  LUT2 id00566 (
    .ADR0(id02404),
    .ADR1(id02401),
    .O(id02408)
  );

  defparam id00567.INIT = 16'h9669;
  LUT4 id00567 (
    .ADR0(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x2 ),
    .O(id02404)
  );

  defparam id00568.INIT = 8'hE8;
  LUT3 id00568 (
    .ADR0(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x2 ),
    .O(id02401)
  );

  defparam id00569.INIT = 8'hB2;
  LUT3 id00569 (
    .ADR0(id02434),
    .ADR1(id02433),
    .ADR2(id02431),
    .O(id02402)
  );

  defparam id00570.INIT = 8'h35;
  LUT3 id00570 (
    .ADR0(id02432),
    .ADR1(id03085),
    .ADR2(id02430),
    .O(id02439)
  );

  defparam id00571.INIT = 4'h4;
  LUT2 id00571 (
    .ADR0(id02429),
    .ADR1(id02428),
    .O(id02438)
  );

  defparam id00572.INIT = 4'h8;
  LUT2 id00572 (
    .ADR0(id02472),
    .ADR1(id02475),
    .O(id02441)
  );

  defparam id00573.INIT = 4'h8;
  LUT2 id00573 (
    .ADR0(id02474),
    .ADR1(id02473),
    .O(id02427)
  );

  defparam id00574.INIT = 4'h8;
  LUT2 id00574 (
    .ADR0(id02484),
    .ADR1(id02483),
    .O(id02426)
  );

  defparam id00575.INIT = 16'h708F;
  LUT4 id00575 (
    .ADR0(id02424),
    .ADR1(id02425),
    .ADR2(id02400),
    .ADR3(id02419),
    .O(\net_Buf-pad-result[54] )
  );

  defparam id00576.INIT = 8'h1F;
  LUT3 id00576 (
    .ADR0(id02426),
    .ADR1(id02427),
    .ADR2(id02423),
    .O(id02400)
  );

  defparam id00577.INIT = 4'h6;
  LUT2 id00577 (
    .ADR0(id02416),
    .ADR1(id02418),
    .O(id02419)
  );

  defparam id00578.INIT = 4'h8;
  LUT2 id00578 (
    .ADR0(id02440),
    .ADR1(id02441),
    .O(id02416)
  );

  defparam id00579.INIT = 8'h1E;
  LUT3 id00579 (
    .ADR0(id02417),
    .ADR1(id02420),
    .ADR2(id02409),
    .O(id02418)
  );

  defparam id00580.INIT = 4'h8;
  LUT2 id00580 (
    .ADR0(id02436),
    .ADR1(id02438),
    .O(id02417)
  );

  defparam id00581.INIT = 4'h4;
  LUT2 id00581 (
    .ADR0(id02439),
    .ADR1(id02435),
    .O(id02420)
  );

  defparam id00582.INIT = 4'h9;
  LUT2 id00582 (
    .ADR0(id02410),
    .ADR1(id02413),
    .O(id02409)
  );

  defparam id00583.INIT = 8'h35;
  LUT3 id00583 (
    .ADR0(id02407),
    .ADR1(id02402),
    .ADR2(id02437),
    .O(id02410)
  );

  defparam id00584.INIT = 4'h6;
  LUT2 id00584 (
    .ADR0(id02415),
    .ADR1(id02414),
    .O(id02413)
  );

  defparam id00585.INIT = 16'h9669;
  LUT4 id00585 (
    .ADR0(id02412),
    .ADR1(id02411),
    .ADR2(id02456),
    .ADR3(id02455),
    .O(id02415)
  );

  defparam id00586.INIT = 8'h35;
  LUT3 id00586 (
    .ADR0(id02401),
    .ADR1(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x0 ),
    .ADR2(id02404),
    .O(id02412)
  );

  defparam id00587.INIT = 4'h9;
  LUT2 id00587 (
    .ADR0(id02457),
    .ADR1(id02459),
    .O(id02411)
  );

  defparam id00588.INIT = 16'h9669;
  LUT4 id00588 (
    .ADR0(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x2 ),
    .O(id02457)
  );

  defparam id00589.INIT = 8'hE8;
  LUT3 id00589 (
    .ADR0(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x2 ),
    .O(id02459)
  );

  defparam id00590.INIT = 16'h6000;
  LUT4 id00590 (
    .ADR0(\u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 ),
    .O(id02456)
  );

  defparam id00591.INIT = 8'h78;
  LUT3 id00591 (
    .ADR0(\u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[40].u_compressor42_cell.x3 ),
    .O(id02455)
  );

  defparam id00592.INIT = 8'hB2;
  LUT3 id00592 (
    .ADR0(id02405),
    .ADR1(id02406),
    .ADR2(id02408),
    .O(id02414)
  );

  defparam id00593.INIT = 8'h1E;
  LUT3 id00593 (
    .ADR0(id02452),
    .ADR1(id02460),
    .ADR2(id02458),
    .O(\net_Buf-pad-result[55] )
  );

  defparam id00594.INIT = 16'h8F00;
  LUT4 id00594 (
    .ADR0(id02425),
    .ADR1(id02424),
    .ADR2(id02400),
    .ADR3(id02419),
    .O(id02452)
  );

  defparam id00595.INIT = 4'h8;
  LUT2 id00595 (
    .ADR0(id02416),
    .ADR1(id02418),
    .O(id02460)
  );

  defparam id00596.INIT = 4'h6;
  LUT2 id00596 (
    .ADR0(id02453),
    .ADR1(id02454),
    .O(id02458)
  );

  defparam id00597.INIT = 4'h8;
  LUT2 id00597 (
    .ADR0(id02417),
    .ADR1(id02409),
    .O(id02453)
  );

  defparam id00598.INIT = 4'h6;
  LUT2 id00598 (
    .ADR0(id02471),
    .ADR1(id02468),
    .O(id02454)
  );

  defparam id00599.INIT = 4'h8;
  LUT2 id00599 (
    .ADR0(id02420),
    .ADR1(id02409),
    .O(id02471)
  );

  defparam id00600.INIT = 4'h6;
  LUT2 id00600 (
    .ADR0(id02467),
    .ADR1(id02470),
    .O(id02468)
  );

  defparam id00601.INIT = 4'h4;
  LUT2 id00601 (
    .ADR0(id02410),
    .ADR1(id02413),
    .O(id02467)
  );

  defparam id00602.INIT = 4'h9;
  LUT2 id00602 (
    .ADR0(id02469),
    .ADR1(id03177),
    .O(id02470)
  );

  defparam id00603.INIT = 8'h35;
  LUT3 id00603 (
    .ADR0(id02455),
    .ADR1(id02414),
    .ADR2(id02415),
    .O(id02469)
  );

  defparam id00604.INIT = 4'h6;
  LUT2 id00604 (
    .ADR0(id03157),
    .ADR1(id03160),
    .O(id03177)
  );

  defparam id00605.INIT = 16'h9669;
  LUT4 id00605 (
    .ADR0(id03159),
    .ADR1(id02462),
    .ADR2(id02461),
    .ADR3(VCC_NET),
    .O(id03157)
  );

  defparam id00606.INIT = 8'h35;
  LUT3 id00606 (
    .ADR0(id02459),
    .ADR1(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x0 ),
    .ADR2(id02457),
    .O(id03159)
  );

  defparam id00607.INIT = 4'h9;
  LUT2 id00607 (
    .ADR0(id02463),
    .ADR1(id02466),
    .O(id02462)
  );

  defparam id00608.INIT = 16'h9669;
  LUT4 id00608 (
    .ADR0(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x2 ),
    .O(id02463)
  );

  defparam id00609.INIT = 8'hE8;
  LUT3 id00609 (
    .ADR0(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x2 ),
    .O(id02466)
  );

  defparam id00610.INIT = 8'h80;
  LUT3 id00610 (
    .ADR0(\u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[40].u_compressor42_cell.x3 ),
    .O(id02461)
  );

  defparam id00611.INIT = 8'hD4;
  LUT3 id00611 (
    .ADR0(id02412),
    .ADR1(id02411),
    .ADR2(id02456),
    .O(id03160)
  );

  defparam id00612.INIT = 16'h708F;
  LUT4 id00612 (
    .ADR0(id02452),
    .ADR1(id02458),
    .ADR2(id02465),
    .ADR3(id02464),
    .O(\net_Buf-pad-result[56] )
  );

  defparam id00613.INIT = 8'h17;
  LUT3 id00613 (
    .ADR0(id02460),
    .ADR1(id02453),
    .ADR2(id02454),
    .O(id02465)
  );

  defparam id00614.INIT = 4'h6;
  LUT2 id00614 (
    .ADR0(id02693),
    .ADR1(id02692),
    .O(id02464)
  );

  defparam id00615.INIT = 4'h8;
  LUT2 id00615 (
    .ADR0(id02471),
    .ADR1(id02468),
    .O(id02693)
  );

  defparam id00616.INIT = 8'h1E;
  LUT3 id00616 (
    .ADR0(id02696),
    .ADR1(id02698),
    .ADR2(id02699),
    .O(id02692)
  );

  defparam id00617.INIT = 4'h8;
  LUT2 id00617 (
    .ADR0(id02467),
    .ADR1(id02470),
    .O(id02696)
  );

  defparam id00618.INIT = 4'h4;
  LUT2 id00618 (
    .ADR0(id02469),
    .ADR1(id03177),
    .O(id02698)
  );

  defparam id00619.INIT = 4'h9;
  LUT2 id00619 (
    .ADR0(id02697),
    .ADR1(id02694),
    .O(id02699)
  );

  defparam id00620.INIT = 8'h35;
  LUT3 id00620 (
    .ADR0(VCC_NET),
    .ADR1(id03160),
    .ADR2(id03157),
    .O(id02697)
  );

  defparam id00621.INIT = 4'h6;
  LUT2 id00621 (
    .ADR0(id02695),
    .ADR1(id02708),
    .O(id02694)
  );

  defparam id00622.INIT = 16'h53AC;
  LUT4 id00622 (
    .ADR0(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x0 ),
    .ADR1(id02466),
    .ADR2(id02463),
    .ADR3(id02709),
    .O(id02695)
  );

  defparam id00623.INIT = 4'h9;
  LUT2 id00623 (
    .ADR0(id02707),
    .ADR1(id02710),
    .O(id02709)
  );

  defparam id00624.INIT = 16'h9669;
  LUT4 id00624 (
    .ADR0(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x2 ),
    .O(id02707)
  );

  defparam id00625.INIT = 8'hE8;
  LUT3 id00625 (
    .ADR0(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x2 ),
    .O(id02710)
  );

  defparam id00626.INIT = 8'hD4;
  LUT3 id00626 (
    .ADR0(id03159),
    .ADR1(id02462),
    .ADR2(id02461),
    .O(id02708)
  );

  defparam id00627.INIT = 16'hE11E;
  LUT4 id00627 (
    .ADR0(id02706),
    .ADR1(id02705),
    .ADR2(id02688),
    .ADR3(id02690),
    .O(\net_Buf-pad-result[57] )
  );

  defparam id00628.INIT = 16'h8F00;
  LUT4 id00628 (
    .ADR0(id02452),
    .ADR1(id02458),
    .ADR2(id02465),
    .ADR3(id02464),
    .O(id02706)
  );

  defparam id00629.INIT = 4'h8;
  LUT2 id00629 (
    .ADR0(id02693),
    .ADR1(id02692),
    .O(id02705)
  );

  defparam id00630.INIT = 4'h8;
  LUT2 id00630 (
    .ADR0(id02696),
    .ADR1(id02699),
    .O(id02688)
  );

  defparam id00631.INIT = 8'h1E;
  LUT3 id00631 (
    .ADR0(id02687),
    .ADR1(id02691),
    .ADR2(id02689),
    .O(id02690)
  );

  defparam id00632.INIT = 4'h8;
  LUT2 id00632 (
    .ADR0(id02698),
    .ADR1(id02699),
    .O(id02687)
  );

  defparam id00633.INIT = 4'h4;
  LUT2 id00633 (
    .ADR0(id02697),
    .ADR1(id02694),
    .O(id02691)
  );

  defparam id00634.INIT = 4'h6;
  LUT2 id00634 (
    .ADR0(id02686),
    .ADR1(id02703),
    .O(id02689)
  );

  defparam id00635.INIT = 4'h8;
  LUT2 id00635 (
    .ADR0(id02695),
    .ADR1(id02708),
    .O(id02686)
  );

  defparam id00636.INIT = 4'h6;
  LUT2 id00636 (
    .ADR0(id02684),
    .ADR1(id02683),
    .O(id02703)
  );

  defparam id00637.INIT = 16'hCA00;
  LUT4 id00637 (
    .ADR0(id02466),
    .ADR1(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x0 ),
    .ADR2(id02463),
    .ADR3(id02709),
    .O(id02684)
  );

  defparam id00638.INIT = 16'h53AC;
  LUT4 id00638 (
    .ADR0(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x0 ),
    .ADR1(id02710),
    .ADR2(id02707),
    .ADR3(id02685),
    .O(id02683)
  );

  defparam id00639.INIT = 4'h9;
  LUT2 id00639 (
    .ADR0(id02780),
    .ADR1(id02782),
    .O(id02685)
  );

  defparam id00640.INIT = 16'h9669;
  LUT4 id00640 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x2 ),
    .O(id02780)
  );

  defparam id00641.INIT = 8'hE8;
  LUT3 id00641 (
    .ADR0(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x2 ),
    .O(id02782)
  );

  defparam id00642.INIT = 8'h69;
  LUT3 id00642 (
    .ADR0(id02783),
    .ADR1(id02781),
    .ADR2(id02779),
    .O(\net_Buf-pad-result[58] )
  );

  defparam id00643.INIT = 16'h1117;
  LUT4 id00643 (
    .ADR0(id02688),
    .ADR1(id02690),
    .ADR2(id02706),
    .ADR3(id02705),
    .O(id02783)
  );

  defparam id00644.INIT = 4'h8;
  LUT2 id00644 (
    .ADR0(id02687),
    .ADR1(id02689),
    .O(id02781)
  );

  defparam id00645.INIT = 4'h9;
  LUT2 id00645 (
    .ADR0(id02772),
    .ADR1(id02778),
    .O(id02779)
  );

  defparam id00646.INIT = 4'h8;
  LUT2 id00646 (
    .ADR0(id02691),
    .ADR1(id02689),
    .O(id02772)
  );

  defparam id00647.INIT = 8'hE1;
  LUT3 id00647 (
    .ADR0(id02775),
    .ADR1(id02777),
    .ADR2(id02776),
    .O(id02778)
  );

  defparam id00648.INIT = 4'h8;
  LUT2 id00648 (
    .ADR0(id02686),
    .ADR1(id02703),
    .O(id02775)
  );

  defparam id00649.INIT = 4'h8;
  LUT2 id00649 (
    .ADR0(id02684),
    .ADR1(id02683),
    .O(id02777)
  );

  defparam id00650.INIT = 4'h6;
  LUT2 id00650 (
    .ADR0(id02774),
    .ADR1(id02773),
    .O(id02776)
  );

  defparam id00651.INIT = 16'hCA00;
  LUT4 id00651 (
    .ADR0(id02710),
    .ADR1(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x0 ),
    .ADR2(id02707),
    .ADR3(id02685),
    .O(id02774)
  );

  defparam id00652.INIT = 16'h53AC;
  LUT4 id00652 (
    .ADR0(VCC_NET),
    .ADR1(id02782),
    .ADR2(id02780),
    .ADR3(id02758),
    .O(id02773)
  );

  defparam id00653.INIT = 16'h17E8;
  LUT4 id00653 (
    .ADR0(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id02760),
    .O(id02758)
  );

  defparam id00654.INIT = 8'h96;
  LUT3 id00654 (
    .ADR0(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x2 ),
    .O(id02760)
  );

  defparam id00655.INIT = 16'h2BD4;
  LUT4 id00655 (
    .ADR0(id02783),
    .ADR1(id02781),
    .ADR2(id02779),
    .ADR3(id02761),
    .O(\net_Buf-pad-result[59] )
  );

  defparam id00656.INIT = 4'h6;
  LUT2 id00656 (
    .ADR0(id02759),
    .ADR1(id02762),
    .O(id02761)
  );

  defparam id00657.INIT = 4'h4;
  LUT2 id00657 (
    .ADR0(id02778),
    .ADR1(id02772),
    .O(id02759)
  );

  defparam id00658.INIT = 4'h6;
  LUT2 id00658 (
    .ADR0(id02763),
    .ADR1(id02769),
    .O(id02762)
  );

  defparam id00659.INIT = 4'h8;
  LUT2 id00659 (
    .ADR0(id02775),
    .ADR1(id02776),
    .O(id02763)
  );

  defparam id00660.INIT = 8'h1E;
  LUT3 id00660 (
    .ADR0(id02770),
    .ADR1(id02768),
    .ADR2(id02771),
    .O(id02769)
  );

  defparam id00661.INIT = 4'h8;
  LUT2 id00661 (
    .ADR0(id02777),
    .ADR1(id02776),
    .O(id02770)
  );

  defparam id00662.INIT = 4'h8;
  LUT2 id00662 (
    .ADR0(id02774),
    .ADR1(id02773),
    .O(id02768)
  );

  defparam id00663.INIT = 4'h6;
  LUT2 id00663 (
    .ADR0(id02767),
    .ADR1(id02766),
    .O(id02771)
  );

  defparam id00664.INIT = 16'hCA00;
  LUT4 id00664 (
    .ADR0(id02782),
    .ADR1(VCC_NET),
    .ADR2(id02780),
    .ADR3(id02758),
    .O(id02767)
  );

  defparam id00665.INIT = 4'h6;
  LUT2 id00665 (
    .ADR0(id02444),
    .ADR1(id02446),
    .O(id02766)
  );

  defparam id00666.INIT = 16'hE800;
  LUT4 id00666 (
    .ADR0(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x2 ),
    .ADR3(id02760),
    .O(id02444)
  );

  defparam id00667.INIT = 16'h6996;
  LUT4 id00667 (
    .ADR0(id02447),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x2 ),
    .O(id02446)
  );

  defparam id00668.INIT = 8'hE8;
  LUT3 id00668 (
    .ADR0(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x2 ),
    .O(id02447)
  );

  defparam id00669.INIT = 8'h1E;
  LUT3 id00669 (
    .ADR0(id02445),
    .ADR1(id02765),
    .ADR2(id02764),
    .O(\net_Buf-pad-result[60] )
  );

  defparam id00670.INIT = 16'hD400;
  LUT4 id00670 (
    .ADR0(id02783),
    .ADR1(id02781),
    .ADR2(id02779),
    .ADR3(id02761),
    .O(id02445)
  );

  defparam id00671.INIT = 4'h8;
  LUT2 id00671 (
    .ADR0(id02759),
    .ADR1(id02762),
    .O(id02765)
  );

  defparam id00672.INIT = 8'h1E;
  LUT3 id00672 (
    .ADR0(id02517),
    .ADR1(id02519),
    .ADR2(id02520),
    .O(id02764)
  );

  defparam id00673.INIT = 4'h8;
  LUT2 id00673 (
    .ADR0(id02763),
    .ADR1(id02769),
    .O(id02517)
  );

  defparam id00674.INIT = 4'h8;
  LUT2 id00674 (
    .ADR0(id02770),
    .ADR1(id02771),
    .O(id02519)
  );

  defparam id00675.INIT = 4'h6;
  LUT2 id00675 (
    .ADR0(id02518),
    .ADR1(id02516),
    .O(id02520)
  );

  defparam id00676.INIT = 4'h8;
  LUT2 id00676 (
    .ADR0(id02768),
    .ADR1(id02771),
    .O(id02518)
  );

  defparam id00677.INIT = 8'h69;
  LUT3 id00677 (
    .ADR0(id02515),
    .ADR1(id02593),
    .ADR2(id02594),
    .O(id02516)
  );

  defparam id00678.INIT = 4'h8;
  LUT2 id00678 (
    .ADR0(id02767),
    .ADR1(id02766),
    .O(id02515)
  );

  defparam id00679.INIT = 4'h1;
  LUT2 id00679 (
    .ADR0(id02592),
    .ADR1(id02591),
    .O(id02593)
  );

  defparam id00680.INIT = 4'h8;
  LUT2 id00680 (
    .ADR0(id02444),
    .ADR1(id02446),
    .O(id02592)
  );

  defparam id00681.INIT = 16'h9600;
  LUT4 id00681 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x2 ),
    .ADR3(id02447),
    .O(id02591)
  );

  defparam id00682.INIT = 8'h96;
  LUT3 id00682 (
    .ADR0(id02513),
    .ADR1(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ),
    .O(id02594)
  );

  defparam id00683.INIT = 8'hE8;
  LUT3 id00683 (
    .ADR0(VCC_NET),
    .ADR1(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x2 ),
    .O(id02513)
  );

  defparam id00684.INIT = 8'h69;
  LUT3 id00684 (
    .ADR0(id02514),
    .ADR1(id02589),
    .ADR2(id02587),
    .O(\net_Buf-pad-result[61] )
  );

  defparam id00685.INIT = 16'h001F;
  LUT4 id00685 (
    .ADR0(id02765),
    .ADR1(id02445),
    .ADR2(id02764),
    .ADR3(id02588),
    .O(id02514)
  );

  defparam id00686.INIT = 4'h8;
  LUT2 id00686 (
    .ADR0(id02517),
    .ADR1(id02520),
    .O(id02588)
  );

  defparam id00687.INIT = 4'h8;
  LUT2 id00687 (
    .ADR0(id02519),
    .ADR1(id02520),
    .O(id02589)
  );

  defparam id00688.INIT = 4'h6;
  LUT2 id00688 (
    .ADR0(id02590),
    .ADR1(id02586),
    .O(id02587)
  );

  defparam id00689.INIT = 4'h8;
  LUT2 id00689 (
    .ADR0(id02518),
    .ADR1(id02516),
    .O(id02590)
  );

  defparam id00690.INIT = 16'h9669;
  LUT4 id00690 (
    .ADR0(id02585),
    .ADR1(id02596),
    .ADR2(id02597),
    .ADR3(id03717),
    .O(id02586)
  );

  defparam id00691.INIT = 4'h8;
  LUT2 id00691 (
    .ADR0(id02594),
    .ADR1(id02515),
    .O(id02585)
  );

  defparam id00692.INIT = 4'h8;
  LUT2 id00692 (
    .ADR0(id02592),
    .ADR1(id02594),
    .O(id02596)
  );

  defparam id00693.INIT = 16'h7117;
  LUT4 id00693 (
    .ADR0(id02591),
    .ADR1(id02513),
    .ADR2(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ),
    .O(id02597)
  );

  defparam id00694.INIT = 16'h8778;
  LUT4 id00694 (
    .ADR0(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(\u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 ),
    .ADR3(VCC_NET),
    .O(id03717)
  );

  defparam id00695.INIT = 8'h69;
  LUT3 id00695 (
    .ADR0(id03718),
    .ADR1(id03721),
    .ADR2(id03722),
    .O(\net_Buf-pad-result[62] )
  );

  defparam id00696.INIT = 8'h2B;
  LUT3 id00696 (
    .ADR0(id02514),
    .ADR1(id02589),
    .ADR2(id02587),
    .O(id03718)
  );

  defparam id00697.INIT = 4'h8;
  LUT2 id00697 (
    .ADR0(id02590),
    .ADR1(id02586),
    .O(id03721)
  );

  defparam id00698.INIT = 8'h94;
  LUT3 id00698 (
    .ADR0(id03723),
    .ADR1(id03725),
    .ADR2(id03726),
    .O(id03722)
  );

  defparam id00699.INIT = 8'h1F;
  LUT3 id00699 (
    .ADR0(id02585),
    .ADR1(id02596),
    .ADR2(id03717),
    .O(id03725)
  );

  defparam id00700.INIT = 8'h80;
  LUT3 id00700 (
    .ADR0(id02591),
    .ADR1(id02594),
    .ADR2(id03717),
    .O(id03723)
  );

  defparam id00701.INIT = 4'h9;
  LUT2 id00701 (
    .ADR0(id03724),
    .ADR1(id03720),
    .O(id03726)
  );

  defparam id00702.INIT = 16'h6000;
  LUT4 id00702 (
    .ADR0(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ),
    .ADR1(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ),
    .ADR2(id02513),
    .ADR3(id03717),
    .O(id03724)
  );

  defparam id00703.INIT = 16'h07F8;
  LUT4 id00703 (
    .ADR0(\u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(id03719),
    .ADR3(\u_compressor42_l0_3.CELLS[40].u_compressor42_cell.x3 ),
    .O(id03720)
  );

  defparam id00704.INIT = 16'h6000;
  LUT4 id00704 (
    .ADR0(\u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 ),
    .O(id03719)
  );

  defparam id00705.INIT = 16'h2BD4;
  LUT4 id00705 (
    .ADR0(id03718),
    .ADR1(id03721),
    .ADR2(id03722),
    .ADR3(id03714),
    .O(\net_Buf-pad-result[63] )
  );

  defparam id00706.INIT = 8'h96;
  LUT3 id00706 (
    .ADR0(id03715),
    .ADR1(id03713),
    .ADR2(id03716),
    .O(id03714)
  );

  defparam id00707.INIT = 8'hB2;
  LUT3 id00707 (
    .ADR0(id03725),
    .ADR1(id03723),
    .ADR2(id03726),
    .O(id03715)
  );

  defparam id00708.INIT = 8'hD3;
  LUT3 id00708 (
    .ADR0(id03724),
    .ADR1(id03719),
    .ADR2(id03720),
    .O(id03713)
  );

  defparam id00709.INIT = 16'h7F80;
  LUT4 id00709 (
    .ADR0(\u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 ),
    .ADR1(VCC_NET),
    .ADR2(\u_compressor42_l0_3.CELLS[40].u_compressor42_cell.x3 ),
    .ADR3(VCC_NET),
    .O(id03716)
  );

  defparam id00710.INIT = 8'h69;
  LUT3 id00710 (
    .ADR0(id03895),
    .ADR1(id03901),
    .ADR2(id03896),
    .O(\net_Buf-pad-result[4] )
  );

  defparam id00711.INIT = 4'h1;
  LUT2 id00711 (
    .ADR0(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 ),
    .O(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x0 )
  );

  defparam id00712.INIT = 8'h70;
  LUT3 id00712 (
    .ADR0(\net_Buf-pad-multiplier[8] ),
    .ADR1(\net_Buf-pad-multiplier[7] ),
    .ADR2(\net_Buf-pad-multiplier[9] ),
    .O(\DECODE_GEN[4].u_booth_enc.partial_reverse )
  );

  defparam id00713.INIT = 8'h70;
  LUT3 id00713 (
    .ADR0(\net_Buf-pad-multiplier[10] ),
    .ADR1(\net_Buf-pad-multiplier[9] ),
    .ADR2(\net_Buf-pad-multiplier[11] ),
    .O(\DECODE_GEN[5].u_booth_enc.partial_reverse )
  );

  defparam id00714.INIT = 8'h70;
  LUT3 id00714 (
    .ADR0(\net_Buf-pad-multiplier[12] ),
    .ADR1(\net_Buf-pad-multiplier[11] ),
    .ADR2(\net_Buf-pad-multiplier[13] ),
    .O(\DECODE_GEN[6].u_booth_enc.partial_reverse )
  );

  defparam id00715.INIT = 8'h70;
  LUT3 id00715 (
    .ADR0(\net_Buf-pad-multiplier[14] ),
    .ADR1(\net_Buf-pad-multiplier[13] ),
    .ADR2(\net_Buf-pad-multiplier[15] ),
    .O(\DECODE_GEN[7].u_booth_enc.partial_reverse )
  );

  defparam id00716.INIT = 8'h70;
  LUT3 id00716 (
    .ADR0(\net_Buf-pad-multiplier[16] ),
    .ADR1(\net_Buf-pad-multiplier[15] ),
    .ADR2(\net_Buf-pad-multiplier[17] ),
    .O(\DECODE_GEN[8].u_booth_enc.partial_reverse )
  );

  defparam id00717.INIT = 8'h70;
  LUT3 id00717 (
    .ADR0(\net_Buf-pad-multiplier[18] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplier[19] ),
    .O(\DECODE_GEN[9].u_booth_enc.partial_reverse )
  );

  defparam id00718.INIT = 8'h70;
  LUT3 id00718 (
    .ADR0(\net_Buf-pad-multiplier[20] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplier[21] ),
    .O(\DECODE_GEN[10].u_booth_enc.partial_reverse )
  );

  defparam id00719.INIT = 8'h70;
  LUT3 id00719 (
    .ADR0(\net_Buf-pad-multiplier[22] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplier[23] ),
    .O(\DECODE_GEN[11].u_booth_enc.partial_reverse )
  );

  defparam id00720.INIT = 8'h70;
  LUT3 id00720 (
    .ADR0(\net_Buf-pad-multiplier[24] ),
    .ADR1(\net_Buf-pad-multiplier[23] ),
    .ADR2(\net_Buf-pad-multiplier[25] ),
    .O(\DECODE_GEN[12].u_booth_enc.partial_reverse )
  );

  defparam id00721.INIT = 8'h70;
  LUT3 id00721 (
    .ADR0(\net_Buf-pad-multiplier[26] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplier[27] ),
    .O(\DECODE_GEN[13].u_booth_enc.partial_reverse )
  );

  defparam id00722.INIT = 8'h70;
  LUT3 id00722 (
    .ADR0(\net_Buf-pad-multiplier[28] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplier[29] ),
    .O(\DECODE_GEN[14].u_booth_enc.partial_reverse )
  );

  defparam id00723.INIT = 8'h70;
  LUT3 id00723 (
    .ADR0(\net_Buf-pad-multiplier[2] ),
    .ADR1(\net_Buf-pad-multiplier[1] ),
    .ADR2(\net_Buf-pad-multiplier[3] ),
    .O(\DECODE_GEN[1].u_booth_enc.partial_reverse )
  );

  defparam id00724.INIT = 8'h70;
  LUT3 id00724 (
    .ADR0(\net_Buf-pad-multiplier[4] ),
    .ADR1(\net_Buf-pad-multiplier[3] ),
    .ADR2(\net_Buf-pad-multiplier[5] ),
    .O(\DECODE_GEN[2].u_booth_enc.partial_reverse )
  );

  defparam id00725.INIT = 8'h70;
  LUT3 id00725 (
    .ADR0(\net_Buf-pad-multiplier[6] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplier[7] ),
    .O(\DECODE_GEN[3].u_booth_enc.partial_reverse )
  );

  defparam id00726.INIT = 16'h0305;
  LUT4 id00726 (
    .ADR0(id04327),
    .ADR1(id04328),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x3 )
  );

  defparam id00727.INIT = 4'h9;
  LUT2 id00727 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[7] ),
    .O(id04328)
  );

  defparam id00728.INIT = 4'h9;
  LUT2 id00728 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[6] ),
    .O(id04327)
  );

  defparam id00729.INIT = 8'h81;
  LUT3 id00729 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplier[6] ),
    .O(id04321)
  );

  defparam id00730.INIT = 4'h6;
  LUT2 id00730 (
    .ADR0(\net_Buf-pad-multiplier[5] ),
    .ADR1(\net_Buf-pad-multiplier[6] ),
    .O(id04322)
  );

  defparam id00731.INIT = 16'h0503;
  LUT4 id00731 (
    .ADR0(id04319),
    .ADR1(id04328),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x3 )
  );

  defparam id00732.INIT = 4'h9;
  LUT2 id00732 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[8] ),
    .O(id04319)
  );

  defparam id00733.INIT = 16'h0503;
  LUT4 id00733 (
    .ADR0(id04320),
    .ADR1(id04319),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x3 )
  );

  defparam id00734.INIT = 4'h9;
  LUT2 id00734 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[9] ),
    .O(id04320)
  );

  defparam id00735.INIT = 16'h0503;
  LUT4 id00735 (
    .ADR0(id04325),
    .ADR1(id04320),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x3 )
  );

  defparam id00736.INIT = 4'h9;
  LUT2 id00736 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[10] ),
    .O(id04325)
  );

  defparam id00737.INIT = 16'h0503;
  LUT4 id00737 (
    .ADR0(id04326),
    .ADR1(id04325),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x3 )
  );

  defparam id00738.INIT = 4'h9;
  LUT2 id00738 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[11] ),
    .O(id04326)
  );

  defparam id00739.INIT = 16'h0503;
  LUT4 id00739 (
    .ADR0(id04323),
    .ADR1(id04326),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x3 )
  );

  defparam id00740.INIT = 4'h9;
  LUT2 id00740 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[12] ),
    .O(id04323)
  );

  defparam id00741.INIT = 16'h0503;
  LUT4 id00741 (
    .ADR0(id04324),
    .ADR1(id04323),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x3 )
  );

  defparam id00742.INIT = 4'h9;
  LUT2 id00742 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[13] ),
    .O(id04324)
  );

  defparam id00743.INIT = 16'h0503;
  LUT4 id00743 (
    .ADR0(id04313),
    .ADR1(id04324),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x3 )
  );

  defparam id00744.INIT = 4'h9;
  LUT2 id00744 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[14] ),
    .O(id04313)
  );

  defparam id00745.INIT = 16'h0503;
  LUT4 id00745 (
    .ADR0(id04314),
    .ADR1(id04313),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x3 )
  );

  defparam id00746.INIT = 4'h9;
  LUT2 id00746 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[15] ),
    .O(id04314)
  );

  defparam id00747.INIT = 16'h0503;
  LUT4 id00747 (
    .ADR0(id04311),
    .ADR1(id04314),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x3 )
  );

  defparam id00748.INIT = 4'h9;
  LUT2 id00748 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[16] ),
    .O(id04311)
  );

  defparam id00749.INIT = 16'h0503;
  LUT4 id00749 (
    .ADR0(id04312),
    .ADR1(id04311),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x3 )
  );

  defparam id00750.INIT = 4'h9;
  LUT2 id00750 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[17] ),
    .O(id04312)
  );

  defparam id00751.INIT = 16'h0503;
  LUT4 id00751 (
    .ADR0(id04317),
    .ADR1(id04312),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x3 )
  );

  defparam id00752.INIT = 4'h9;
  LUT2 id00752 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[18] ),
    .O(id04317)
  );

  defparam id00753.INIT = 16'h0503;
  LUT4 id00753 (
    .ADR0(id04318),
    .ADR1(id04317),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x3 )
  );

  defparam id00754.INIT = 4'h9;
  LUT2 id00754 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[19] ),
    .O(id04318)
  );

  defparam id00755.INIT = 16'h0503;
  LUT4 id00755 (
    .ADR0(id04315),
    .ADR1(id04318),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x3 )
  );

  defparam id00756.INIT = 4'h9;
  LUT2 id00756 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[20] ),
    .O(id04315)
  );

  defparam id00757.INIT = 16'h0503;
  LUT4 id00757 (
    .ADR0(id04316),
    .ADR1(id04315),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x3 )
  );

  defparam id00758.INIT = 4'h9;
  LUT2 id00758 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[21] ),
    .O(id04316)
  );

  defparam id00759.INIT = 16'h0503;
  LUT4 id00759 (
    .ADR0(id04305),
    .ADR1(id04316),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x3 )
  );

  defparam id00760.INIT = 4'h9;
  LUT2 id00760 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[22] ),
    .O(id04305)
  );

  defparam id00761.INIT = 16'h0503;
  LUT4 id00761 (
    .ADR0(id04306),
    .ADR1(id04305),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x3 )
  );

  defparam id00762.INIT = 4'h9;
  LUT2 id00762 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[23] ),
    .O(id04306)
  );

  defparam id00763.INIT = 16'h0503;
  LUT4 id00763 (
    .ADR0(id04303),
    .ADR1(id04306),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x3 )
  );

  defparam id00764.INIT = 4'h9;
  LUT2 id00764 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[24] ),
    .O(id04303)
  );

  defparam id00765.INIT = 16'h0503;
  LUT4 id00765 (
    .ADR0(id04304),
    .ADR1(id04303),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x3 )
  );

  defparam id00766.INIT = 4'h9;
  LUT2 id00766 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[25] ),
    .O(id04304)
  );

  defparam id00767.INIT = 16'h0503;
  LUT4 id00767 (
    .ADR0(id04309),
    .ADR1(id04304),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x3 )
  );

  defparam id00768.INIT = 4'h9;
  LUT2 id00768 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[26] ),
    .O(id04309)
  );

  defparam id00769.INIT = 16'h0503;
  LUT4 id00769 (
    .ADR0(id04310),
    .ADR1(id04309),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x3 )
  );

  defparam id00770.INIT = 4'h9;
  LUT2 id00770 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[27] ),
    .O(id04310)
  );

  defparam id00771.INIT = 16'h0503;
  LUT4 id00771 (
    .ADR0(id04307),
    .ADR1(id04310),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x3 )
  );

  defparam id00772.INIT = 4'h9;
  LUT2 id00772 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[28] ),
    .O(id04307)
  );

  defparam id00773.INIT = 16'h0503;
  LUT4 id00773 (
    .ADR0(id04308),
    .ADR1(id04307),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x3 )
  );

  defparam id00774.INIT = 4'h9;
  LUT2 id00774 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[29] ),
    .O(id04308)
  );

  defparam id00775.INIT = 16'h0503;
  LUT4 id00775 (
    .ADR0(id04355),
    .ADR1(id04308),
    .ADR2(id04321),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x3 )
  );

  defparam id00776.INIT = 4'h9;
  LUT2 id00776 (
    .ADR0(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR1(\net_Buf-pad-multiplicand[30] ),
    .O(id04355)
  );

  defparam id00777.INIT = 16'h3307;
  LUT4 id00777 (
    .ADR0(id04321),
    .ADR1(\u_compressor42_l0_0.CELLS[38].u_compressor42_cell.x3 ),
    .ADR2(id04355),
    .ADR3(id04322),
    .O(\u_compressor42_l0_0.CELLS[37].u_compressor42_cell.x3 )
  );

  defparam id00778.INIT = 8'hEB;
  LUT3 id00778 (
    .ADR0(id04321),
    .ADR1(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_0.CELLS[38].u_compressor42_cell.x3 )
  );

  defparam id00779.INIT = 16'h1760;
  LUT4 id00779 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(\u_compressor42_l0_1.CELLS[2].u_compressor42_cell.x0 )
  );

  defparam id00780.INIT = 16'h00BE;
  LUT4 id00780 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04353),
    .O(\u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 )
  );

  defparam id00781.INIT = 4'h6;
  LUT2 id00781 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .O(id04356)
  );

  defparam id00782.INIT = 16'hE817;
  LUT4 id00782 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04353)
  );

  defparam id00783.INIT = 16'h00BE;
  LUT4 id00783 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04354),
    .O(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x0 )
  );

  defparam id00784.INIT = 16'hE817;
  LUT4 id00784 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04354)
  );

  defparam id00785.INIT = 16'h00BE;
  LUT4 id00785 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04359),
    .O(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x0 )
  );

  defparam id00786.INIT = 16'hE817;
  LUT4 id00786 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04359)
  );

  defparam id00787.INIT = 16'h00BE;
  LUT4 id00787 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04360),
    .O(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x0 )
  );

  defparam id00788.INIT = 16'hE817;
  LUT4 id00788 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04360)
  );

  defparam id00789.INIT = 16'h00BE;
  LUT4 id00789 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04357),
    .O(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x0 )
  );

  defparam id00790.INIT = 16'hE817;
  LUT4 id00790 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04357)
  );

  defparam id00791.INIT = 16'h00BE;
  LUT4 id00791 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04358),
    .O(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x0 )
  );

  defparam id00792.INIT = 16'hE817;
  LUT4 id00792 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04358)
  );

  defparam id00793.INIT = 16'h00BE;
  LUT4 id00793 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04347),
    .O(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x0 )
  );

  defparam id00794.INIT = 16'hE817;
  LUT4 id00794 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04347)
  );

  defparam id00795.INIT = 16'h00BE;
  LUT4 id00795 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04348),
    .O(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x0 )
  );

  defparam id00796.INIT = 16'hE817;
  LUT4 id00796 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04348)
  );

  defparam id00797.INIT = 16'h00BE;
  LUT4 id00797 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04345),
    .O(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x0 )
  );

  defparam id00798.INIT = 16'hE817;
  LUT4 id00798 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04345)
  );

  defparam id00799.INIT = 16'h00BE;
  LUT4 id00799 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04346),
    .O(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x0 )
  );

  defparam id00800.INIT = 16'hE817;
  LUT4 id00800 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04346)
  );

  defparam id00801.INIT = 16'h00BE;
  LUT4 id00801 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04351),
    .O(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x0 )
  );

  defparam id00802.INIT = 16'hE817;
  LUT4 id00802 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04351)
  );

  defparam id00803.INIT = 16'h00BE;
  LUT4 id00803 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04352),
    .O(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x0 )
  );

  defparam id00804.INIT = 16'hE817;
  LUT4 id00804 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04352)
  );

  defparam id00805.INIT = 16'h00BE;
  LUT4 id00805 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04349),
    .O(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x0 )
  );

  defparam id00806.INIT = 16'hE817;
  LUT4 id00806 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04349)
  );

  defparam id00807.INIT = 16'h00BE;
  LUT4 id00807 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04350),
    .O(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x0 )
  );

  defparam id00808.INIT = 16'hE817;
  LUT4 id00808 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04350)
  );

  defparam id00809.INIT = 16'h00BE;
  LUT4 id00809 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04339),
    .O(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x0 )
  );

  defparam id00810.INIT = 16'hE817;
  LUT4 id00810 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04339)
  );

  defparam id00811.INIT = 16'h00BE;
  LUT4 id00811 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id04340),
    .O(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x0 )
  );

  defparam id00812.INIT = 16'hE817;
  LUT4 id00812 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04340)
  );

  defparam id00813.INIT = 16'h00BE;
  LUT4 id00813 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04337),
    .O(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x0 )
  );

  defparam id00814.INIT = 16'hE817;
  LUT4 id00814 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04337)
  );

  defparam id00815.INIT = 16'h00BE;
  LUT4 id00815 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04338),
    .O(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x0 )
  );

  defparam id00816.INIT = 16'hE817;
  LUT4 id00816 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04338)
  );

  defparam id00817.INIT = 16'h00BE;
  LUT4 id00817 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04343),
    .O(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x0 )
  );

  defparam id00818.INIT = 16'hE817;
  LUT4 id00818 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04343)
  );

  defparam id00819.INIT = 16'h00BE;
  LUT4 id00819 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04344),
    .O(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x0 )
  );

  defparam id00820.INIT = 16'hE817;
  LUT4 id00820 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04344)
  );

  defparam id00821.INIT = 16'h00BE;
  LUT4 id00821 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04341),
    .O(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x0 )
  );

  defparam id00822.INIT = 16'hE817;
  LUT4 id00822 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04341)
  );

  defparam id00823.INIT = 16'h00BE;
  LUT4 id00823 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04342),
    .O(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x0 )
  );

  defparam id00824.INIT = 16'hE817;
  LUT4 id00824 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04342)
  );

  defparam id00825.INIT = 16'h00BE;
  LUT4 id00825 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04331),
    .O(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x0 )
  );

  defparam id00826.INIT = 16'hE817;
  LUT4 id00826 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04331)
  );

  defparam id00827.INIT = 16'h00BE;
  LUT4 id00827 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04332),
    .O(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x0 )
  );

  defparam id00828.INIT = 16'hE817;
  LUT4 id00828 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04332)
  );

  defparam id00829.INIT = 16'h00BE;
  LUT4 id00829 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04329),
    .O(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x0 )
  );

  defparam id00830.INIT = 16'hE817;
  LUT4 id00830 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04329)
  );

  defparam id00831.INIT = 16'h00BE;
  LUT4 id00831 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04330),
    .O(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x0 )
  );

  defparam id00832.INIT = 16'hE817;
  LUT4 id00832 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04330)
  );

  defparam id00833.INIT = 16'h00BE;
  LUT4 id00833 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04335),
    .O(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x0 )
  );

  defparam id00834.INIT = 16'hE817;
  LUT4 id00834 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04335)
  );

  defparam id00835.INIT = 16'h00BE;
  LUT4 id00835 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04336),
    .O(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x0 )
  );

  defparam id00836.INIT = 16'hE817;
  LUT4 id00836 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04336)
  );

  defparam id00837.INIT = 16'h00BE;
  LUT4 id00837 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04333),
    .O(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x0 )
  );

  defparam id00838.INIT = 16'hE817;
  LUT4 id00838 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04333)
  );

  defparam id00839.INIT = 16'h00BE;
  LUT4 id00839 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04334),
    .O(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x0 )
  );

  defparam id00840.INIT = 16'hE817;
  LUT4 id00840 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04334)
  );

  defparam id00841.INIT = 16'h00BE;
  LUT4 id00841 (
    .ADR0(id04356),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04265),
    .O(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x0 )
  );

  defparam id00842.INIT = 16'hE817;
  LUT4 id00842 (
    .ADR0(\net_Buf-pad-multiplier[7] ),
    .ADR1(\net_Buf-pad-multiplier[8] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[9] ),
    .O(id04265)
  );

  defparam id00843.INIT = 16'hABD5;
  LUT4 id00843 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[7] ),
    .ADR2(\net_Buf-pad-multiplier[8] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x0 )
  );

  defparam id00844.INIT = 16'h1760;
  LUT4 id00844 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 )
  );

  defparam id00845.INIT = 16'h00BE;
  LUT4 id00845 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04263),
    .O(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 )
  );

  defparam id00846.INIT = 4'h6;
  LUT2 id00846 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .O(id04266)
  );

  defparam id00847.INIT = 16'hE817;
  LUT4 id00847 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04263)
  );

  defparam id00848.INIT = 16'h00BE;
  LUT4 id00848 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04264),
    .O(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x1 )
  );

  defparam id00849.INIT = 16'hE817;
  LUT4 id00849 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04264)
  );

  defparam id00850.INIT = 16'h00BE;
  LUT4 id00850 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04269),
    .O(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x1 )
  );

  defparam id00851.INIT = 16'hE817;
  LUT4 id00851 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04269)
  );

  defparam id00852.INIT = 16'h00BE;
  LUT4 id00852 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04270),
    .O(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x1 )
  );

  defparam id00853.INIT = 16'hE817;
  LUT4 id00853 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04270)
  );

  defparam id00854.INIT = 16'h00BE;
  LUT4 id00854 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04267),
    .O(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x1 )
  );

  defparam id00855.INIT = 16'hE817;
  LUT4 id00855 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04267)
  );

  defparam id00856.INIT = 16'h00BE;
  LUT4 id00856 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04268),
    .O(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x1 )
  );

  defparam id00857.INIT = 16'hE817;
  LUT4 id00857 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04268)
  );

  defparam id00858.INIT = 16'h00BE;
  LUT4 id00858 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04257),
    .O(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x1 )
  );

  defparam id00859.INIT = 16'hE817;
  LUT4 id00859 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04257)
  );

  defparam id00860.INIT = 16'h00BE;
  LUT4 id00860 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04258),
    .O(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x1 )
  );

  defparam id00861.INIT = 16'hE817;
  LUT4 id00861 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04258)
  );

  defparam id00862.INIT = 16'h00BE;
  LUT4 id00862 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04255),
    .O(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x1 )
  );

  defparam id00863.INIT = 16'hE817;
  LUT4 id00863 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04255)
  );

  defparam id00864.INIT = 16'h00BE;
  LUT4 id00864 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04256),
    .O(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x1 )
  );

  defparam id00865.INIT = 16'hE817;
  LUT4 id00865 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04256)
  );

  defparam id00866.INIT = 16'h00BE;
  LUT4 id00866 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04261),
    .O(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x1 )
  );

  defparam id00867.INIT = 16'hE817;
  LUT4 id00867 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04261)
  );

  defparam id00868.INIT = 16'h00BE;
  LUT4 id00868 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04262),
    .O(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x1 )
  );

  defparam id00869.INIT = 16'hE817;
  LUT4 id00869 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04262)
  );

  defparam id00870.INIT = 16'h00BE;
  LUT4 id00870 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04259),
    .O(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x1 )
  );

  defparam id00871.INIT = 16'hE817;
  LUT4 id00871 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04259)
  );

  defparam id00872.INIT = 16'h00BE;
  LUT4 id00872 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04260),
    .O(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x1 )
  );

  defparam id00873.INIT = 16'hE817;
  LUT4 id00873 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04260)
  );

  defparam id00874.INIT = 16'h00BE;
  LUT4 id00874 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04249),
    .O(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x1 )
  );

  defparam id00875.INIT = 16'hE817;
  LUT4 id00875 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04249)
  );

  defparam id00876.INIT = 16'h00BE;
  LUT4 id00876 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id04250),
    .O(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x1 )
  );

  defparam id00877.INIT = 16'hE817;
  LUT4 id00877 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04250)
  );

  defparam id00878.INIT = 16'h00BE;
  LUT4 id00878 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04247),
    .O(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x1 )
  );

  defparam id00879.INIT = 16'hE817;
  LUT4 id00879 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04247)
  );

  defparam id00880.INIT = 16'h00BE;
  LUT4 id00880 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04248),
    .O(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x1 )
  );

  defparam id00881.INIT = 16'hE817;
  LUT4 id00881 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04248)
  );

  defparam id00882.INIT = 16'h00BE;
  LUT4 id00882 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04253),
    .O(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x1 )
  );

  defparam id00883.INIT = 16'hE817;
  LUT4 id00883 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04253)
  );

  defparam id00884.INIT = 16'h00BE;
  LUT4 id00884 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04254),
    .O(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x1 )
  );

  defparam id00885.INIT = 16'hE817;
  LUT4 id00885 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04254)
  );

  defparam id00886.INIT = 16'h00BE;
  LUT4 id00886 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04251),
    .O(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x1 )
  );

  defparam id00887.INIT = 16'hE817;
  LUT4 id00887 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04251)
  );

  defparam id00888.INIT = 16'h00BE;
  LUT4 id00888 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04252),
    .O(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x1 )
  );

  defparam id00889.INIT = 16'hE817;
  LUT4 id00889 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04252)
  );

  defparam id00890.INIT = 16'h00BE;
  LUT4 id00890 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04241),
    .O(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x1 )
  );

  defparam id00891.INIT = 16'hE817;
  LUT4 id00891 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04241)
  );

  defparam id00892.INIT = 16'h00BE;
  LUT4 id00892 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04242),
    .O(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x1 )
  );

  defparam id00893.INIT = 16'hE817;
  LUT4 id00893 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04242)
  );

  defparam id00894.INIT = 16'h00BE;
  LUT4 id00894 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04239),
    .O(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x1 )
  );

  defparam id00895.INIT = 16'hE817;
  LUT4 id00895 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04239)
  );

  defparam id00896.INIT = 16'h00BE;
  LUT4 id00896 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04240),
    .O(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x1 )
  );

  defparam id00897.INIT = 16'hE817;
  LUT4 id00897 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04240)
  );

  defparam id00898.INIT = 16'h00BE;
  LUT4 id00898 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04245),
    .O(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x1 )
  );

  defparam id00899.INIT = 16'hE817;
  LUT4 id00899 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04245)
  );

  defparam id00900.INIT = 16'h00BE;
  LUT4 id00900 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04246),
    .O(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x1 )
  );

  defparam id00901.INIT = 16'hE817;
  LUT4 id00901 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04246)
  );

  defparam id00902.INIT = 16'h00BE;
  LUT4 id00902 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04243),
    .O(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x1 )
  );

  defparam id00903.INIT = 16'hE817;
  LUT4 id00903 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04243)
  );

  defparam id00904.INIT = 16'h00BE;
  LUT4 id00904 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04244),
    .O(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x1 )
  );

  defparam id00905.INIT = 16'hE817;
  LUT4 id00905 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04244)
  );

  defparam id00906.INIT = 16'h00BE;
  LUT4 id00906 (
    .ADR0(id04266),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04297),
    .O(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x1 )
  );

  defparam id00907.INIT = 16'hE817;
  LUT4 id00907 (
    .ADR0(\net_Buf-pad-multiplier[9] ),
    .ADR1(\net_Buf-pad-multiplier[10] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[11] ),
    .O(id04297)
  );

  defparam id00908.INIT = 16'hABD5;
  LUT4 id00908 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[9] ),
    .ADR2(\net_Buf-pad-multiplier[10] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x1 )
  );

  defparam id00909.INIT = 16'h1760;
  LUT4 id00909 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x2 )
  );

  defparam id00910.INIT = 16'h00BE;
  LUT4 id00910 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04295),
    .O(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x2 )
  );

  defparam id00911.INIT = 4'h6;
  LUT2 id00911 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .O(id04298)
  );

  defparam id00912.INIT = 16'hE817;
  LUT4 id00912 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04295)
  );

  defparam id00913.INIT = 16'h00BE;
  LUT4 id00913 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04296),
    .O(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x2 )
  );

  defparam id00914.INIT = 16'hE817;
  LUT4 id00914 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04296)
  );

  defparam id00915.INIT = 16'h00BE;
  LUT4 id00915 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04301),
    .O(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x2 )
  );

  defparam id00916.INIT = 16'hE817;
  LUT4 id00916 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04301)
  );

  defparam id00917.INIT = 16'h00BE;
  LUT4 id00917 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04302),
    .O(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x2 )
  );

  defparam id00918.INIT = 16'hE817;
  LUT4 id00918 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04302)
  );

  defparam id00919.INIT = 16'h00BE;
  LUT4 id00919 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04299),
    .O(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x2 )
  );

  defparam id00920.INIT = 16'hE817;
  LUT4 id00920 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04299)
  );

  defparam id00921.INIT = 16'h00BE;
  LUT4 id00921 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04300),
    .O(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x2 )
  );

  defparam id00922.INIT = 16'hE817;
  LUT4 id00922 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04300)
  );

  defparam id00923.INIT = 16'h00BE;
  LUT4 id00923 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04289),
    .O(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x2 )
  );

  defparam id00924.INIT = 16'hE817;
  LUT4 id00924 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04289)
  );

  defparam id00925.INIT = 16'h00BE;
  LUT4 id00925 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04290),
    .O(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x2 )
  );

  defparam id00926.INIT = 16'hE817;
  LUT4 id00926 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04290)
  );

  defparam id00927.INIT = 16'h00BE;
  LUT4 id00927 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04287),
    .O(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x2 )
  );

  defparam id00928.INIT = 16'hE817;
  LUT4 id00928 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04287)
  );

  defparam id00929.INIT = 16'h00BE;
  LUT4 id00929 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04288),
    .O(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x2 )
  );

  defparam id00930.INIT = 16'hE817;
  LUT4 id00930 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04288)
  );

  defparam id00931.INIT = 16'h00BE;
  LUT4 id00931 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04293),
    .O(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x2 )
  );

  defparam id00932.INIT = 16'hE817;
  LUT4 id00932 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04293)
  );

  defparam id00933.INIT = 16'h00BE;
  LUT4 id00933 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04294),
    .O(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x2 )
  );

  defparam id00934.INIT = 16'hE817;
  LUT4 id00934 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04294)
  );

  defparam id00935.INIT = 16'h00BE;
  LUT4 id00935 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04291),
    .O(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x2 )
  );

  defparam id00936.INIT = 16'hE817;
  LUT4 id00936 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04291)
  );

  defparam id00937.INIT = 16'h00BE;
  LUT4 id00937 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04292),
    .O(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x2 )
  );

  defparam id00938.INIT = 16'hE817;
  LUT4 id00938 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04292)
  );

  defparam id00939.INIT = 16'h00BE;
  LUT4 id00939 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04281),
    .O(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x2 )
  );

  defparam id00940.INIT = 16'hE817;
  LUT4 id00940 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04281)
  );

  defparam id00941.INIT = 16'h00BE;
  LUT4 id00941 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id04282),
    .O(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x2 )
  );

  defparam id00942.INIT = 16'hE817;
  LUT4 id00942 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04282)
  );

  defparam id00943.INIT = 16'h00BE;
  LUT4 id00943 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04279),
    .O(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x2 )
  );

  defparam id00944.INIT = 16'hE817;
  LUT4 id00944 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04279)
  );

  defparam id00945.INIT = 16'h00BE;
  LUT4 id00945 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04280),
    .O(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x2 )
  );

  defparam id00946.INIT = 16'hE817;
  LUT4 id00946 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04280)
  );

  defparam id00947.INIT = 16'h00BE;
  LUT4 id00947 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04285),
    .O(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x2 )
  );

  defparam id00948.INIT = 16'hE817;
  LUT4 id00948 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04285)
  );

  defparam id00949.INIT = 16'h00BE;
  LUT4 id00949 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04286),
    .O(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x2 )
  );

  defparam id00950.INIT = 16'hE817;
  LUT4 id00950 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04286)
  );

  defparam id00951.INIT = 16'h00BE;
  LUT4 id00951 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04283),
    .O(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x2 )
  );

  defparam id00952.INIT = 16'hE817;
  LUT4 id00952 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04283)
  );

  defparam id00953.INIT = 16'h00BE;
  LUT4 id00953 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04284),
    .O(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x2 )
  );

  defparam id00954.INIT = 16'hE817;
  LUT4 id00954 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04284)
  );

  defparam id00955.INIT = 16'h00BE;
  LUT4 id00955 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04273),
    .O(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x2 )
  );

  defparam id00956.INIT = 16'hE817;
  LUT4 id00956 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04273)
  );

  defparam id00957.INIT = 16'h00BE;
  LUT4 id00957 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04274),
    .O(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x2 )
  );

  defparam id00958.INIT = 16'hE817;
  LUT4 id00958 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04274)
  );

  defparam id00959.INIT = 16'h00BE;
  LUT4 id00959 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04271),
    .O(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x2 )
  );

  defparam id00960.INIT = 16'hE817;
  LUT4 id00960 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04271)
  );

  defparam id00961.INIT = 16'h00BE;
  LUT4 id00961 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04272),
    .O(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x2 )
  );

  defparam id00962.INIT = 16'hE817;
  LUT4 id00962 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04272)
  );

  defparam id00963.INIT = 16'h00BE;
  LUT4 id00963 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04277),
    .O(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x2 )
  );

  defparam id00964.INIT = 16'hE817;
  LUT4 id00964 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04277)
  );

  defparam id00965.INIT = 16'h00BE;
  LUT4 id00965 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04278),
    .O(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x2 )
  );

  defparam id00966.INIT = 16'hE817;
  LUT4 id00966 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04278)
  );

  defparam id00967.INIT = 16'h00BE;
  LUT4 id00967 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04275),
    .O(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x2 )
  );

  defparam id00968.INIT = 16'hE817;
  LUT4 id00968 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04275)
  );

  defparam id00969.INIT = 16'h00BE;
  LUT4 id00969 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04276),
    .O(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x2 )
  );

  defparam id00970.INIT = 16'hE817;
  LUT4 id00970 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04276)
  );

  defparam id00971.INIT = 16'h00BE;
  LUT4 id00971 (
    .ADR0(id04298),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04451),
    .O(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x2 )
  );

  defparam id00972.INIT = 16'hE817;
  LUT4 id00972 (
    .ADR0(\net_Buf-pad-multiplier[11] ),
    .ADR1(\net_Buf-pad-multiplier[12] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[13] ),
    .O(id04451)
  );

  defparam id00973.INIT = 16'hABD5;
  LUT4 id00973 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[11] ),
    .ADR2(\net_Buf-pad-multiplier[12] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x2 )
  );

  defparam id00974.INIT = 16'h1760;
  LUT4 id00974 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x3 )
  );

  defparam id00975.INIT = 16'h00BE;
  LUT4 id00975 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04449),
    .O(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x3 )
  );

  defparam id00976.INIT = 4'h6;
  LUT2 id00976 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .O(id04452)
  );

  defparam id00977.INIT = 16'hE817;
  LUT4 id00977 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04449)
  );

  defparam id00978.INIT = 16'h00BE;
  LUT4 id00978 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04450),
    .O(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x3 )
  );

  defparam id00979.INIT = 16'hE817;
  LUT4 id00979 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04450)
  );

  defparam id00980.INIT = 16'h00BE;
  LUT4 id00980 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04455),
    .O(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x3 )
  );

  defparam id00981.INIT = 16'hE817;
  LUT4 id00981 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04455)
  );

  defparam id00982.INIT = 16'h00BE;
  LUT4 id00982 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04456),
    .O(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x3 )
  );

  defparam id00983.INIT = 16'hE817;
  LUT4 id00983 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04456)
  );

  defparam id00984.INIT = 16'h00BE;
  LUT4 id00984 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04453),
    .O(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x3 )
  );

  defparam id00985.INIT = 16'hE817;
  LUT4 id00985 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04453)
  );

  defparam id00986.INIT = 16'h00BE;
  LUT4 id00986 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04454),
    .O(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x3 )
  );

  defparam id00987.INIT = 16'hE817;
  LUT4 id00987 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04454)
  );

  defparam id00988.INIT = 16'h00BE;
  LUT4 id00988 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04443),
    .O(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x3 )
  );

  defparam id00989.INIT = 16'hE817;
  LUT4 id00989 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04443)
  );

  defparam id00990.INIT = 16'h00BE;
  LUT4 id00990 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04444),
    .O(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x3 )
  );

  defparam id00991.INIT = 16'hE817;
  LUT4 id00991 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04444)
  );

  defparam id00992.INIT = 16'h00BE;
  LUT4 id00992 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04441),
    .O(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x3 )
  );

  defparam id00993.INIT = 16'hE817;
  LUT4 id00993 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04441)
  );

  defparam id00994.INIT = 16'h00BE;
  LUT4 id00994 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04442),
    .O(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x3 )
  );

  defparam id00995.INIT = 16'hE817;
  LUT4 id00995 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04442)
  );

  defparam id00996.INIT = 16'h00BE;
  LUT4 id00996 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04447),
    .O(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x3 )
  );

  defparam id00997.INIT = 16'hE817;
  LUT4 id00997 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04447)
  );

  defparam id00998.INIT = 16'h00BE;
  LUT4 id00998 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04448),
    .O(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x3 )
  );

  defparam id00999.INIT = 16'hE817;
  LUT4 id00999 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04448)
  );

  defparam id01000.INIT = 16'h00BE;
  LUT4 id01000 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04445),
    .O(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x3 )
  );

  defparam id01001.INIT = 16'hE817;
  LUT4 id01001 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04445)
  );

  defparam id01002.INIT = 16'h00BE;
  LUT4 id01002 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04446),
    .O(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x3 )
  );

  defparam id01003.INIT = 16'hE817;
  LUT4 id01003 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04446)
  );

  defparam id01004.INIT = 16'h00BE;
  LUT4 id01004 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04435),
    .O(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x3 )
  );

  defparam id01005.INIT = 16'hE817;
  LUT4 id01005 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04435)
  );

  defparam id01006.INIT = 16'h00BE;
  LUT4 id01006 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id04436),
    .O(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x3 )
  );

  defparam id01007.INIT = 16'hE817;
  LUT4 id01007 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04436)
  );

  defparam id01008.INIT = 16'h00BE;
  LUT4 id01008 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04433),
    .O(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x3 )
  );

  defparam id01009.INIT = 16'hE817;
  LUT4 id01009 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04433)
  );

  defparam id01010.INIT = 16'h00BE;
  LUT4 id01010 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04434),
    .O(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x3 )
  );

  defparam id01011.INIT = 16'hE817;
  LUT4 id01011 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04434)
  );

  defparam id01012.INIT = 16'h00BE;
  LUT4 id01012 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04439),
    .O(\u_compressor42_l0_1.CELLS[27].u_compressor42_cell.x3 )
  );

  defparam id01013.INIT = 16'hE817;
  LUT4 id01013 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04439)
  );

  defparam id01014.INIT = 16'h00BE;
  LUT4 id01014 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04440),
    .O(\u_compressor42_l0_1.CELLS[28].u_compressor42_cell.x3 )
  );

  defparam id01015.INIT = 16'hE817;
  LUT4 id01015 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04440)
  );

  defparam id01016.INIT = 16'h00BE;
  LUT4 id01016 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04437),
    .O(\u_compressor42_l0_1.CELLS[29].u_compressor42_cell.x3 )
  );

  defparam id01017.INIT = 16'hE817;
  LUT4 id01017 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04437)
  );

  defparam id01018.INIT = 16'h00BE;
  LUT4 id01018 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04438),
    .O(\u_compressor42_l0_1.CELLS[30].u_compressor42_cell.x3 )
  );

  defparam id01019.INIT = 16'hE817;
  LUT4 id01019 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04438)
  );

  defparam id01020.INIT = 16'h00BE;
  LUT4 id01020 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04427),
    .O(\u_compressor42_l0_1.CELLS[31].u_compressor42_cell.x3 )
  );

  defparam id01021.INIT = 16'hE817;
  LUT4 id01021 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04427)
  );

  defparam id01022.INIT = 16'h00BE;
  LUT4 id01022 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04428),
    .O(\u_compressor42_l0_1.CELLS[32].u_compressor42_cell.x3 )
  );

  defparam id01023.INIT = 16'hE817;
  LUT4 id01023 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04428)
  );

  defparam id01024.INIT = 16'h00BE;
  LUT4 id01024 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04425),
    .O(\u_compressor42_l0_1.CELLS[33].u_compressor42_cell.x3 )
  );

  defparam id01025.INIT = 16'hE817;
  LUT4 id01025 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04425)
  );

  defparam id01026.INIT = 16'h00BE;
  LUT4 id01026 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04426),
    .O(\u_compressor42_l0_1.CELLS[34].u_compressor42_cell.x3 )
  );

  defparam id01027.INIT = 16'hE817;
  LUT4 id01027 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04426)
  );

  defparam id01028.INIT = 16'h00BE;
  LUT4 id01028 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04431),
    .O(\u_compressor42_l0_1.CELLS[35].u_compressor42_cell.x3 )
  );

  defparam id01029.INIT = 16'hE817;
  LUT4 id01029 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04431)
  );

  defparam id01030.INIT = 16'h00BE;
  LUT4 id01030 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04432),
    .O(\u_compressor42_l0_1.CELLS[36].u_compressor42_cell.x3 )
  );

  defparam id01031.INIT = 16'hE817;
  LUT4 id01031 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04432)
  );

  defparam id01032.INIT = 16'h00BE;
  LUT4 id01032 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04429),
    .O(\u_compressor42_l0_1.CELLS[37].u_compressor42_cell.x3 )
  );

  defparam id01033.INIT = 16'hE817;
  LUT4 id01033 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04429)
  );

  defparam id01034.INIT = 16'h00BE;
  LUT4 id01034 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04430),
    .O(\u_compressor42_l0_1.CELLS[38].u_compressor42_cell.x3 )
  );

  defparam id01035.INIT = 16'hE817;
  LUT4 id01035 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04430)
  );

  defparam id01036.INIT = 16'h00BE;
  LUT4 id01036 (
    .ADR0(id04452),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04483),
    .O(\u_compressor42_l0_1.CELLS[39].u_compressor42_cell.x3 )
  );

  defparam id01037.INIT = 16'hE817;
  LUT4 id01037 (
    .ADR0(\net_Buf-pad-multiplier[13] ),
    .ADR1(\net_Buf-pad-multiplier[14] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[15] ),
    .O(id04483)
  );

  defparam id01038.INIT = 16'hABD5;
  LUT4 id01038 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[13] ),
    .ADR2(\net_Buf-pad-multiplier[14] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_1.CELLS[40].u_compressor42_cell.x3 )
  );

  defparam id01039.INIT = 16'h1760;
  LUT4 id01039 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(\u_compressor42_l0_2.CELLS[2].u_compressor42_cell.x0 )
  );

  defparam id01040.INIT = 16'h7D00;
  LUT4 id01040 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04481),
    .O(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 )
  );

  defparam id01041.INIT = 4'h6;
  LUT2 id01041 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .O(id04484)
  );

  defparam id01042.INIT = 16'h75AE;
  LUT4 id01042 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04481)
  );

  defparam id01043.INIT = 16'h00BE;
  LUT4 id01043 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04482),
    .O(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x0 )
  );

  defparam id01044.INIT = 16'hE817;
  LUT4 id01044 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04482)
  );

  defparam id01045.INIT = 16'h7D00;
  LUT4 id01045 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04487),
    .O(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x0 )
  );

  defparam id01046.INIT = 16'h75AE;
  LUT4 id01046 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04487)
  );

  defparam id01047.INIT = 16'h7D00;
  LUT4 id01047 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04488),
    .O(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x0 )
  );

  defparam id01048.INIT = 16'h75AE;
  LUT4 id01048 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04488)
  );

  defparam id01049.INIT = 16'h7D00;
  LUT4 id01049 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04485),
    .O(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x0 )
  );

  defparam id01050.INIT = 16'h75AE;
  LUT4 id01050 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04485)
  );

  defparam id01051.INIT = 16'h7D00;
  LUT4 id01051 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04486),
    .O(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x0 )
  );

  defparam id01052.INIT = 16'h75AE;
  LUT4 id01052 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04486)
  );

  defparam id01053.INIT = 16'h7D00;
  LUT4 id01053 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04475),
    .O(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x0 )
  );

  defparam id01054.INIT = 16'h75AE;
  LUT4 id01054 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04475)
  );

  defparam id01055.INIT = 16'h7D00;
  LUT4 id01055 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04476),
    .O(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x0 )
  );

  defparam id01056.INIT = 16'h75AE;
  LUT4 id01056 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04476)
  );

  defparam id01057.INIT = 16'h00BE;
  LUT4 id01057 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04473),
    .O(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x0 )
  );

  defparam id01058.INIT = 16'hE817;
  LUT4 id01058 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04473)
  );

  defparam id01059.INIT = 16'h7D00;
  LUT4 id01059 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04474),
    .O(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x0 )
  );

  defparam id01060.INIT = 16'h75AE;
  LUT4 id01060 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04474)
  );

  defparam id01061.INIT = 16'h00BE;
  LUT4 id01061 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04479),
    .O(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x0 )
  );

  defparam id01062.INIT = 16'hE817;
  LUT4 id01062 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04479)
  );

  defparam id01063.INIT = 16'h00BE;
  LUT4 id01063 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04480),
    .O(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x0 )
  );

  defparam id01064.INIT = 16'hE817;
  LUT4 id01064 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04480)
  );

  defparam id01065.INIT = 16'h00BE;
  LUT4 id01065 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04477),
    .O(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x0 )
  );

  defparam id01066.INIT = 16'hE817;
  LUT4 id01066 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04477)
  );

  defparam id01067.INIT = 16'h7D00;
  LUT4 id01067 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04478),
    .O(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x0 )
  );

  defparam id01068.INIT = 16'h75AE;
  LUT4 id01068 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04478)
  );

  defparam id01069.INIT = 16'h00BE;
  LUT4 id01069 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04467),
    .O(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x0 )
  );

  defparam id01070.INIT = 16'hE817;
  LUT4 id01070 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04467)
  );

  defparam id01071.INIT = 16'h7D00;
  LUT4 id01071 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04468),
    .O(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x0 )
  );

  defparam id01072.INIT = 16'h75AE;
  LUT4 id01072 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04468)
  );

  defparam id01073.INIT = 16'h7D00;
  LUT4 id01073 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04465),
    .O(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x0 )
  );

  defparam id01074.INIT = 16'h75AE;
  LUT4 id01074 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04465)
  );

  defparam id01075.INIT = 16'h7D00;
  LUT4 id01075 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04466),
    .O(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x0 )
  );

  defparam id01076.INIT = 16'h75AE;
  LUT4 id01076 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04466)
  );

  defparam id01077.INIT = 16'h7D00;
  LUT4 id01077 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04471),
    .O(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x0 )
  );

  defparam id01078.INIT = 16'h75AE;
  LUT4 id01078 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04471)
  );

  defparam id01079.INIT = 16'h7D00;
  LUT4 id01079 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04472),
    .O(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x0 )
  );

  defparam id01080.INIT = 16'h75AE;
  LUT4 id01080 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04472)
  );

  defparam id01081.INIT = 16'h7D00;
  LUT4 id01081 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04469),
    .O(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x0 )
  );

  defparam id01082.INIT = 16'h75AE;
  LUT4 id01082 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04469)
  );

  defparam id01083.INIT = 16'h7D00;
  LUT4 id01083 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04470),
    .O(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x0 )
  );

  defparam id01084.INIT = 16'h75AE;
  LUT4 id01084 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04470)
  );

  defparam id01085.INIT = 16'h7D00;
  LUT4 id01085 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04459),
    .O(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x0 )
  );

  defparam id01086.INIT = 16'h75AE;
  LUT4 id01086 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04459)
  );

  defparam id01087.INIT = 16'h00BE;
  LUT4 id01087 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04460),
    .O(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x0 )
  );

  defparam id01088.INIT = 16'hE817;
  LUT4 id01088 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04460)
  );

  defparam id01089.INIT = 16'h7D00;
  LUT4 id01089 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04457),
    .O(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x0 )
  );

  defparam id01090.INIT = 16'h75AE;
  LUT4 id01090 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04457)
  );

  defparam id01091.INIT = 16'h00BE;
  LUT4 id01091 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04458),
    .O(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x0 )
  );

  defparam id01092.INIT = 16'hE817;
  LUT4 id01092 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04458)
  );

  defparam id01093.INIT = 16'h7D00;
  LUT4 id01093 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04463),
    .O(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x0 )
  );

  defparam id01094.INIT = 16'h75AE;
  LUT4 id01094 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04463)
  );

  defparam id01095.INIT = 16'h00BE;
  LUT4 id01095 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id04464),
    .O(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x0 )
  );

  defparam id01096.INIT = 16'hE817;
  LUT4 id01096 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04464)
  );

  defparam id01097.INIT = 16'h00BE;
  LUT4 id01097 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04461),
    .O(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x0 )
  );

  defparam id01098.INIT = 16'hE817;
  LUT4 id01098 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04461)
  );

  defparam id01099.INIT = 16'h7D00;
  LUT4 id01099 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04462),
    .O(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x0 )
  );

  defparam id01100.INIT = 16'h75AE;
  LUT4 id01100 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[16] ),
    .O(id04462)
  );

  defparam id01101.INIT = 16'h00BE;
  LUT4 id01101 (
    .ADR0(id04484),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04387),
    .O(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x0 )
  );

  defparam id01102.INIT = 16'hE817;
  LUT4 id01102 (
    .ADR0(\net_Buf-pad-multiplier[15] ),
    .ADR1(\net_Buf-pad-multiplier[16] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[17] ),
    .O(id04387)
  );

  defparam id01103.INIT = 16'hABD5;
  LUT4 id01103 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[15] ),
    .ADR2(\net_Buf-pad-multiplier[16] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x0 )
  );

  defparam id01104.INIT = 16'h1760;
  LUT4 id01104 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x1 )
  );

  defparam id01105.INIT = 16'h00BE;
  LUT4 id01105 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04385),
    .O(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 )
  );

  defparam id01106.INIT = 4'h6;
  LUT2 id01106 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .O(id04388)
  );

  defparam id01107.INIT = 16'hE817;
  LUT4 id01107 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04385)
  );

  defparam id01108.INIT = 16'h00BE;
  LUT4 id01108 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id04386),
    .O(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x1 )
  );

  defparam id01109.INIT = 16'hE817;
  LUT4 id01109 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04386)
  );

  defparam id01110.INIT = 16'h00BE;
  LUT4 id01110 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04391),
    .O(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x1 )
  );

  defparam id01111.INIT = 16'hE817;
  LUT4 id01111 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04391)
  );

  defparam id01112.INIT = 16'h7D00;
  LUT4 id01112 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id04392),
    .O(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x1 )
  );

  defparam id01113.INIT = 16'h75AE;
  LUT4 id01113 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04392)
  );

  defparam id01114.INIT = 16'h7D00;
  LUT4 id01114 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04389),
    .O(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x1 )
  );

  defparam id01115.INIT = 16'h75AE;
  LUT4 id01115 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04389)
  );

  defparam id01116.INIT = 16'h7D00;
  LUT4 id01116 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04390),
    .O(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x1 )
  );

  defparam id01117.INIT = 16'h75AE;
  LUT4 id01117 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04390)
  );

  defparam id01118.INIT = 16'h7D00;
  LUT4 id01118 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04379),
    .O(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x1 )
  );

  defparam id01119.INIT = 16'h75AE;
  LUT4 id01119 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04379)
  );

  defparam id01120.INIT = 16'h7D00;
  LUT4 id01120 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id04380),
    .O(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x1 )
  );

  defparam id01121.INIT = 16'h75AE;
  LUT4 id01121 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04380)
  );

  defparam id01122.INIT = 16'h7D00;
  LUT4 id01122 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04377),
    .O(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x1 )
  );

  defparam id01123.INIT = 16'h75AE;
  LUT4 id01123 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04377)
  );

  defparam id01124.INIT = 16'h7D00;
  LUT4 id01124 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04378),
    .O(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x1 )
  );

  defparam id01125.INIT = 16'h75AE;
  LUT4 id01125 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04378)
  );

  defparam id01126.INIT = 16'h00BE;
  LUT4 id01126 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id04383),
    .O(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x1 )
  );

  defparam id01127.INIT = 16'hE817;
  LUT4 id01127 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04383)
  );

  defparam id01128.INIT = 16'h7D00;
  LUT4 id01128 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04384),
    .O(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x1 )
  );

  defparam id01129.INIT = 16'h75AE;
  LUT4 id01129 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04384)
  );

  defparam id01130.INIT = 16'h7D00;
  LUT4 id01130 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04381),
    .O(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x1 )
  );

  defparam id01131.INIT = 16'h75AE;
  LUT4 id01131 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04381)
  );

  defparam id01132.INIT = 16'h7D00;
  LUT4 id01132 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04382),
    .O(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x1 )
  );

  defparam id01133.INIT = 16'h75AE;
  LUT4 id01133 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04382)
  );

  defparam id01134.INIT = 16'h00BE;
  LUT4 id01134 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id04371),
    .O(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x1 )
  );

  defparam id01135.INIT = 16'hE817;
  LUT4 id01135 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04371)
  );

  defparam id01136.INIT = 16'h7D00;
  LUT4 id01136 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04372),
    .O(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x1 )
  );

  defparam id01137.INIT = 16'h75AE;
  LUT4 id01137 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04372)
  );

  defparam id01138.INIT = 16'h7D00;
  LUT4 id01138 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04369),
    .O(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x1 )
  );

  defparam id01139.INIT = 16'h75AE;
  LUT4 id01139 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04369)
  );

  defparam id01140.INIT = 16'h7D00;
  LUT4 id01140 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04370),
    .O(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x1 )
  );

  defparam id01141.INIT = 16'h75AE;
  LUT4 id01141 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04370)
  );

  defparam id01142.INIT = 16'h00BE;
  LUT4 id01142 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id04375),
    .O(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x1 )
  );

  defparam id01143.INIT = 16'hE817;
  LUT4 id01143 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04375)
  );

  defparam id01144.INIT = 16'h7D00;
  LUT4 id01144 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id04376),
    .O(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x1 )
  );

  defparam id01145.INIT = 16'h75AE;
  LUT4 id01145 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04376)
  );

  defparam id01146.INIT = 16'h7D00;
  LUT4 id01146 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04373),
    .O(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x1 )
  );

  defparam id01147.INIT = 16'h75AE;
  LUT4 id01147 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04373)
  );

  defparam id01148.INIT = 16'h7D00;
  LUT4 id01148 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04374),
    .O(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x1 )
  );

  defparam id01149.INIT = 16'h75AE;
  LUT4 id01149 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04374)
  );

  defparam id01150.INIT = 16'h7D00;
  LUT4 id01150 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04363),
    .O(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x1 )
  );

  defparam id01151.INIT = 16'h75AE;
  LUT4 id01151 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04363)
  );

  defparam id01152.INIT = 16'h00BE;
  LUT4 id01152 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04364),
    .O(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x1 )
  );

  defparam id01153.INIT = 16'hE817;
  LUT4 id01153 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04364)
  );

  defparam id01154.INIT = 16'h00BE;
  LUT4 id01154 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04361),
    .O(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x1 )
  );

  defparam id01155.INIT = 16'hE817;
  LUT4 id01155 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04361)
  );

  defparam id01156.INIT = 16'h7D00;
  LUT4 id01156 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04362),
    .O(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x1 )
  );

  defparam id01157.INIT = 16'h75AE;
  LUT4 id01157 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04362)
  );

  defparam id01158.INIT = 16'h00BE;
  LUT4 id01158 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04367),
    .O(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x1 )
  );

  defparam id01159.INIT = 16'hE817;
  LUT4 id01159 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04367)
  );

  defparam id01160.INIT = 16'h7D00;
  LUT4 id01160 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04368),
    .O(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x1 )
  );

  defparam id01161.INIT = 16'h75AE;
  LUT4 id01161 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04368)
  );

  defparam id01162.INIT = 16'h7D00;
  LUT4 id01162 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04365),
    .O(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x1 )
  );

  defparam id01163.INIT = 16'h75AE;
  LUT4 id01163 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04365)
  );

  defparam id01164.INIT = 16'h7D00;
  LUT4 id01164 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04366),
    .O(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x1 )
  );

  defparam id01165.INIT = 16'h75AE;
  LUT4 id01165 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[18] ),
    .O(id04366)
  );

  defparam id01166.INIT = 16'h00BE;
  LUT4 id01166 (
    .ADR0(id04388),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id04419),
    .O(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x1 )
  );

  defparam id01167.INIT = 16'hE817;
  LUT4 id01167 (
    .ADR0(\net_Buf-pad-multiplier[17] ),
    .ADR1(\net_Buf-pad-multiplier[18] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[19] ),
    .O(id04419)
  );

  defparam id01168.INIT = 16'hABD5;
  LUT4 id01168 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[17] ),
    .ADR2(\net_Buf-pad-multiplier[18] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x1 )
  );

  defparam id01169.INIT = 16'h1760;
  LUT4 id01169 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x2 )
  );

  defparam id01170.INIT = 16'h00BE;
  LUT4 id01170 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id04417),
    .O(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x2 )
  );

  defparam id01171.INIT = 4'h6;
  LUT2 id01171 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .O(id04420)
  );

  defparam id01172.INIT = 16'hE817;
  LUT4 id01172 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04417)
  );

  defparam id01173.INIT = 16'h7D00;
  LUT4 id01173 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04418),
    .O(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x2 )
  );

  defparam id01174.INIT = 16'h75AE;
  LUT4 id01174 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04418)
  );

  defparam id01175.INIT = 16'h00BE;
  LUT4 id01175 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id04423),
    .O(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x2 )
  );

  defparam id01176.INIT = 16'hE817;
  LUT4 id01176 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04423)
  );

  defparam id01177.INIT = 16'h00BE;
  LUT4 id01177 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id04424),
    .O(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x2 )
  );

  defparam id01178.INIT = 16'hE817;
  LUT4 id01178 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04424)
  );

  defparam id01179.INIT = 16'h7D00;
  LUT4 id01179 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id04421),
    .O(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x2 )
  );

  defparam id01180.INIT = 16'h75AE;
  LUT4 id01180 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04421)
  );

  defparam id01181.INIT = 16'h7D00;
  LUT4 id01181 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id04422),
    .O(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x2 )
  );

  defparam id01182.INIT = 16'h75AE;
  LUT4 id01182 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04422)
  );

  defparam id01183.INIT = 16'h7D00;
  LUT4 id01183 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04411),
    .O(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x2 )
  );

  defparam id01184.INIT = 16'h75AE;
  LUT4 id01184 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04411)
  );

  defparam id01185.INIT = 16'h00BE;
  LUT4 id01185 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id04412),
    .O(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x2 )
  );

  defparam id01186.INIT = 16'hE817;
  LUT4 id01186 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04412)
  );

  defparam id01187.INIT = 16'h7D00;
  LUT4 id01187 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04409),
    .O(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x2 )
  );

  defparam id01188.INIT = 16'h75AE;
  LUT4 id01188 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04409)
  );

  defparam id01189.INIT = 16'h00BE;
  LUT4 id01189 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id04410),
    .O(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x2 )
  );

  defparam id01190.INIT = 16'hE817;
  LUT4 id01190 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04410)
  );

  defparam id01191.INIT = 16'h7D00;
  LUT4 id01191 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id04415),
    .O(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x2 )
  );

  defparam id01192.INIT = 16'h75AE;
  LUT4 id01192 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04415)
  );

  defparam id01193.INIT = 16'h7D00;
  LUT4 id01193 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04416),
    .O(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x2 )
  );

  defparam id01194.INIT = 16'h75AE;
  LUT4 id01194 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04416)
  );

  defparam id01195.INIT = 16'h00BE;
  LUT4 id01195 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id04413),
    .O(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x2 )
  );

  defparam id01196.INIT = 16'hE817;
  LUT4 id01196 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04413)
  );

  defparam id01197.INIT = 16'h00BE;
  LUT4 id01197 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id04414),
    .O(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x2 )
  );

  defparam id01198.INIT = 16'hE817;
  LUT4 id01198 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04414)
  );

  defparam id01199.INIT = 16'h7D00;
  LUT4 id01199 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id04403),
    .O(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x2 )
  );

  defparam id01200.INIT = 16'h75AE;
  LUT4 id01200 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04403)
  );

  defparam id01201.INIT = 16'h7D00;
  LUT4 id01201 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04404),
    .O(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x2 )
  );

  defparam id01202.INIT = 16'h75AE;
  LUT4 id01202 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04404)
  );

  defparam id01203.INIT = 16'h00BE;
  LUT4 id01203 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id04401),
    .O(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x2 )
  );

  defparam id01204.INIT = 16'hE817;
  LUT4 id01204 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04401)
  );

  defparam id01205.INIT = 16'h00BE;
  LUT4 id01205 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id04402),
    .O(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x2 )
  );

  defparam id01206.INIT = 16'hE817;
  LUT4 id01206 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04402)
  );

  defparam id01207.INIT = 16'h7D00;
  LUT4 id01207 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04407),
    .O(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x2 )
  );

  defparam id01208.INIT = 16'h75AE;
  LUT4 id01208 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04407)
  );

  defparam id01209.INIT = 16'h00BE;
  LUT4 id01209 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id04408),
    .O(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x2 )
  );

  defparam id01210.INIT = 16'hE817;
  LUT4 id01210 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04408)
  );

  defparam id01211.INIT = 16'h7D00;
  LUT4 id01211 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id04405),
    .O(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x2 )
  );

  defparam id01212.INIT = 16'h75AE;
  LUT4 id01212 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04405)
  );

  defparam id01213.INIT = 16'h7D00;
  LUT4 id01213 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id04406),
    .O(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x2 )
  );

  defparam id01214.INIT = 16'h75AE;
  LUT4 id01214 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04406)
  );

  defparam id01215.INIT = 16'h7D00;
  LUT4 id01215 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id04395),
    .O(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x2 )
  );

  defparam id01216.INIT = 16'h75AE;
  LUT4 id01216 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04395)
  );

  defparam id01217.INIT = 16'h7D00;
  LUT4 id01217 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id04396),
    .O(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x2 )
  );

  defparam id01218.INIT = 16'h75AE;
  LUT4 id01218 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04396)
  );

  defparam id01219.INIT = 16'h7D00;
  LUT4 id01219 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04393),
    .O(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x2 )
  );

  defparam id01220.INIT = 16'h75AE;
  LUT4 id01220 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04393)
  );

  defparam id01221.INIT = 16'h00BE;
  LUT4 id01221 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id04394),
    .O(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x2 )
  );

  defparam id01222.INIT = 16'hE817;
  LUT4 id01222 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04394)
  );

  defparam id01223.INIT = 16'h00BE;
  LUT4 id01223 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id04399),
    .O(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x2 )
  );

  defparam id01224.INIT = 16'hE817;
  LUT4 id01224 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04399)
  );

  defparam id01225.INIT = 16'h7D00;
  LUT4 id01225 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id04400),
    .O(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x2 )
  );

  defparam id01226.INIT = 16'h75AE;
  LUT4 id01226 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04400)
  );

  defparam id01227.INIT = 16'h7D00;
  LUT4 id01227 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04397),
    .O(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x2 )
  );

  defparam id01228.INIT = 16'h75AE;
  LUT4 id01228 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[20] ),
    .O(id04397)
  );

  defparam id01229.INIT = 16'h00BE;
  LUT4 id01229 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id04398),
    .O(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x2 )
  );

  defparam id01230.INIT = 16'hE817;
  LUT4 id01230 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id04398)
  );

  defparam id01231.INIT = 16'h00BE;
  LUT4 id01231 (
    .ADR0(id04420),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03817),
    .O(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x2 )
  );

  defparam id01232.INIT = 16'hE817;
  LUT4 id01232 (
    .ADR0(\net_Buf-pad-multiplier[19] ),
    .ADR1(\net_Buf-pad-multiplier[20] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[21] ),
    .O(id03817)
  );

  defparam id01233.INIT = 16'hABD5;
  LUT4 id01233 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[19] ),
    .ADR2(\net_Buf-pad-multiplier[20] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x2 )
  );

  defparam id01234.INIT = 16'h1760;
  LUT4 id01234 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x3 )
  );

  defparam id01235.INIT = 16'h00BE;
  LUT4 id01235 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id03815),
    .O(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x3 )
  );

  defparam id01236.INIT = 4'h6;
  LUT2 id01236 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .O(id03818)
  );

  defparam id01237.INIT = 16'hE817;
  LUT4 id01237 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03815)
  );

  defparam id01238.INIT = 16'h00BE;
  LUT4 id01238 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03816),
    .O(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x3 )
  );

  defparam id01239.INIT = 16'hE817;
  LUT4 id01239 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03816)
  );

  defparam id01240.INIT = 16'h00BE;
  LUT4 id01240 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03821),
    .O(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x3 )
  );

  defparam id01241.INIT = 16'hE817;
  LUT4 id01241 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03821)
  );

  defparam id01242.INIT = 16'h00BE;
  LUT4 id01242 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03822),
    .O(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x3 )
  );

  defparam id01243.INIT = 16'hE817;
  LUT4 id01243 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03822)
  );

  defparam id01244.INIT = 16'h00BE;
  LUT4 id01244 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03819),
    .O(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x3 )
  );

  defparam id01245.INIT = 16'hE817;
  LUT4 id01245 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03819)
  );

  defparam id01246.INIT = 16'h00BE;
  LUT4 id01246 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03820),
    .O(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x3 )
  );

  defparam id01247.INIT = 16'hE817;
  LUT4 id01247 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03820)
  );

  defparam id01248.INIT = 16'h00BE;
  LUT4 id01248 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03809),
    .O(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x3 )
  );

  defparam id01249.INIT = 16'hE817;
  LUT4 id01249 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03809)
  );

  defparam id01250.INIT = 16'h00BE;
  LUT4 id01250 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03810),
    .O(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x3 )
  );

  defparam id01251.INIT = 16'hE817;
  LUT4 id01251 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03810)
  );

  defparam id01252.INIT = 16'h00BE;
  LUT4 id01252 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03807),
    .O(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x3 )
  );

  defparam id01253.INIT = 16'hE817;
  LUT4 id01253 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03807)
  );

  defparam id01254.INIT = 16'h00BE;
  LUT4 id01254 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03808),
    .O(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x3 )
  );

  defparam id01255.INIT = 16'hE817;
  LUT4 id01255 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03808)
  );

  defparam id01256.INIT = 16'h00BE;
  LUT4 id01256 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03813),
    .O(\u_compressor42_l0_2.CELLS[19].u_compressor42_cell.x3 )
  );

  defparam id01257.INIT = 16'hE817;
  LUT4 id01257 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03813)
  );

  defparam id01258.INIT = 16'h00BE;
  LUT4 id01258 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03814),
    .O(\u_compressor42_l0_2.CELLS[20].u_compressor42_cell.x3 )
  );

  defparam id01259.INIT = 16'hE817;
  LUT4 id01259 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03814)
  );

  defparam id01260.INIT = 16'h00BE;
  LUT4 id01260 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03811),
    .O(\u_compressor42_l0_2.CELLS[21].u_compressor42_cell.x3 )
  );

  defparam id01261.INIT = 16'hE817;
  LUT4 id01261 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03811)
  );

  defparam id01262.INIT = 16'h00BE;
  LUT4 id01262 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id03812),
    .O(\u_compressor42_l0_2.CELLS[22].u_compressor42_cell.x3 )
  );

  defparam id01263.INIT = 16'hE817;
  LUT4 id01263 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03812)
  );

  defparam id01264.INIT = 16'h00BE;
  LUT4 id01264 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03801),
    .O(\u_compressor42_l0_2.CELLS[23].u_compressor42_cell.x3 )
  );

  defparam id01265.INIT = 16'hE817;
  LUT4 id01265 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03801)
  );

  defparam id01266.INIT = 16'h00BE;
  LUT4 id01266 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03802),
    .O(\u_compressor42_l0_2.CELLS[24].u_compressor42_cell.x3 )
  );

  defparam id01267.INIT = 16'hE817;
  LUT4 id01267 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03802)
  );

  defparam id01268.INIT = 16'h00BE;
  LUT4 id01268 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03799),
    .O(\u_compressor42_l0_2.CELLS[25].u_compressor42_cell.x3 )
  );

  defparam id01269.INIT = 16'hE817;
  LUT4 id01269 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03799)
  );

  defparam id01270.INIT = 16'h00BE;
  LUT4 id01270 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03800),
    .O(\u_compressor42_l0_2.CELLS[26].u_compressor42_cell.x3 )
  );

  defparam id01271.INIT = 16'hE817;
  LUT4 id01271 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03800)
  );

  defparam id01272.INIT = 16'h00BE;
  LUT4 id01272 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03805),
    .O(\u_compressor42_l0_2.CELLS[27].u_compressor42_cell.x3 )
  );

  defparam id01273.INIT = 16'hE817;
  LUT4 id01273 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03805)
  );

  defparam id01274.INIT = 16'h00BE;
  LUT4 id01274 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03806),
    .O(\u_compressor42_l0_2.CELLS[28].u_compressor42_cell.x3 )
  );

  defparam id01275.INIT = 16'hE817;
  LUT4 id01275 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03806)
  );

  defparam id01276.INIT = 16'h00BE;
  LUT4 id01276 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03803),
    .O(\u_compressor42_l0_2.CELLS[29].u_compressor42_cell.x3 )
  );

  defparam id01277.INIT = 16'hE817;
  LUT4 id01277 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03803)
  );

  defparam id01278.INIT = 16'h00BE;
  LUT4 id01278 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03804),
    .O(\u_compressor42_l0_2.CELLS[30].u_compressor42_cell.x3 )
  );

  defparam id01279.INIT = 16'hE817;
  LUT4 id01279 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03804)
  );

  defparam id01280.INIT = 16'h00BE;
  LUT4 id01280 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03793),
    .O(\u_compressor42_l0_2.CELLS[31].u_compressor42_cell.x3 )
  );

  defparam id01281.INIT = 16'hE817;
  LUT4 id01281 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03793)
  );

  defparam id01282.INIT = 16'h00BE;
  LUT4 id01282 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03794),
    .O(\u_compressor42_l0_2.CELLS[32].u_compressor42_cell.x3 )
  );

  defparam id01283.INIT = 16'hE817;
  LUT4 id01283 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03794)
  );

  defparam id01284.INIT = 16'h00BE;
  LUT4 id01284 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03791),
    .O(\u_compressor42_l0_2.CELLS[33].u_compressor42_cell.x3 )
  );

  defparam id01285.INIT = 16'hE817;
  LUT4 id01285 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03791)
  );

  defparam id01286.INIT = 16'h00BE;
  LUT4 id01286 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03792),
    .O(\u_compressor42_l0_2.CELLS[34].u_compressor42_cell.x3 )
  );

  defparam id01287.INIT = 16'hE817;
  LUT4 id01287 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03792)
  );

  defparam id01288.INIT = 16'h00BE;
  LUT4 id01288 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03797),
    .O(\u_compressor42_l0_2.CELLS[35].u_compressor42_cell.x3 )
  );

  defparam id01289.INIT = 16'hE817;
  LUT4 id01289 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03797)
  );

  defparam id01290.INIT = 16'h00BE;
  LUT4 id01290 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03798),
    .O(\u_compressor42_l0_2.CELLS[36].u_compressor42_cell.x3 )
  );

  defparam id01291.INIT = 16'hE817;
  LUT4 id01291 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03798)
  );

  defparam id01292.INIT = 16'h00BE;
  LUT4 id01292 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03795),
    .O(\u_compressor42_l0_2.CELLS[37].u_compressor42_cell.x3 )
  );

  defparam id01293.INIT = 16'hE817;
  LUT4 id01293 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03795)
  );

  defparam id01294.INIT = 16'h00BE;
  LUT4 id01294 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03796),
    .O(\u_compressor42_l0_2.CELLS[38].u_compressor42_cell.x3 )
  );

  defparam id01295.INIT = 16'hE817;
  LUT4 id01295 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03796)
  );

  defparam id01296.INIT = 16'h00BE;
  LUT4 id01296 (
    .ADR0(id03818),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03849),
    .O(\u_compressor42_l0_2.CELLS[39].u_compressor42_cell.x3 )
  );

  defparam id01297.INIT = 16'hE817;
  LUT4 id01297 (
    .ADR0(\net_Buf-pad-multiplier[21] ),
    .ADR1(\net_Buf-pad-multiplier[22] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[23] ),
    .O(id03849)
  );

  defparam id01298.INIT = 16'hABD5;
  LUT4 id01298 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[21] ),
    .ADR2(\net_Buf-pad-multiplier[22] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_2.CELLS[40].u_compressor42_cell.x3 )
  );

  defparam id01299.INIT = 16'h1760;
  LUT4 id01299 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(\u_compressor42_l0_3.CELLS[2].u_compressor42_cell.x0 )
  );

  defparam id01300.INIT = 16'h7D00;
  LUT4 id01300 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03847),
    .O(\u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 )
  );

  defparam id01301.INIT = 4'h6;
  LUT2 id01301 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .O(id03850)
  );

  defparam id01302.INIT = 16'h75AE;
  LUT4 id01302 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03847)
  );

  defparam id01303.INIT = 16'h7D00;
  LUT4 id01303 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03848),
    .O(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x0 )
  );

  defparam id01304.INIT = 16'h75AE;
  LUT4 id01304 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03848)
  );

  defparam id01305.INIT = 16'h00BE;
  LUT4 id01305 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03853),
    .O(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x0 )
  );

  defparam id01306.INIT = 16'hE817;
  LUT4 id01306 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03853)
  );

  defparam id01307.INIT = 16'h00BE;
  LUT4 id01307 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03854),
    .O(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x0 )
  );

  defparam id01308.INIT = 16'hE817;
  LUT4 id01308 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03854)
  );

  defparam id01309.INIT = 16'h7D00;
  LUT4 id01309 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03851),
    .O(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x0 )
  );

  defparam id01310.INIT = 16'h75AE;
  LUT4 id01310 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03851)
  );

  defparam id01311.INIT = 16'h7D00;
  LUT4 id01311 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03852),
    .O(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x0 )
  );

  defparam id01312.INIT = 16'h75AE;
  LUT4 id01312 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03852)
  );

  defparam id01313.INIT = 16'h7D00;
  LUT4 id01313 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03841),
    .O(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x0 )
  );

  defparam id01314.INIT = 16'h75AE;
  LUT4 id01314 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03841)
  );

  defparam id01315.INIT = 16'h7D00;
  LUT4 id01315 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03842),
    .O(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x0 )
  );

  defparam id01316.INIT = 16'h75AE;
  LUT4 id01316 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03842)
  );

  defparam id01317.INIT = 16'h7D00;
  LUT4 id01317 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03839),
    .O(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x0 )
  );

  defparam id01318.INIT = 16'h75AE;
  LUT4 id01318 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03839)
  );

  defparam id01319.INIT = 16'h00BE;
  LUT4 id01319 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03840),
    .O(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x0 )
  );

  defparam id01320.INIT = 16'hE817;
  LUT4 id01320 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03840)
  );

  defparam id01321.INIT = 16'h7D00;
  LUT4 id01321 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03845),
    .O(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x0 )
  );

  defparam id01322.INIT = 16'h75AE;
  LUT4 id01322 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03845)
  );

  defparam id01323.INIT = 16'h7D00;
  LUT4 id01323 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03846),
    .O(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x0 )
  );

  defparam id01324.INIT = 16'h75AE;
  LUT4 id01324 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03846)
  );

  defparam id01325.INIT = 16'h00BE;
  LUT4 id01325 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03843),
    .O(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x0 )
  );

  defparam id01326.INIT = 16'hE817;
  LUT4 id01326 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03843)
  );

  defparam id01327.INIT = 16'h7D00;
  LUT4 id01327 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03844),
    .O(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x0 )
  );

  defparam id01328.INIT = 16'h75AE;
  LUT4 id01328 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03844)
  );

  defparam id01329.INIT = 16'h7D00;
  LUT4 id01329 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03833),
    .O(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x0 )
  );

  defparam id01330.INIT = 16'h75AE;
  LUT4 id01330 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03833)
  );

  defparam id01331.INIT = 16'h7D00;
  LUT4 id01331 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03834),
    .O(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x0 )
  );

  defparam id01332.INIT = 16'h75AE;
  LUT4 id01332 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03834)
  );

  defparam id01333.INIT = 16'h00BE;
  LUT4 id01333 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03831),
    .O(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x0 )
  );

  defparam id01334.INIT = 16'hE817;
  LUT4 id01334 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03831)
  );

  defparam id01335.INIT = 16'h7D00;
  LUT4 id01335 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03832),
    .O(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x0 )
  );

  defparam id01336.INIT = 16'h75AE;
  LUT4 id01336 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03832)
  );

  defparam id01337.INIT = 16'h7D00;
  LUT4 id01337 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03837),
    .O(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x0 )
  );

  defparam id01338.INIT = 16'h75AE;
  LUT4 id01338 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03837)
  );

  defparam id01339.INIT = 16'h7D00;
  LUT4 id01339 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03838),
    .O(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x0 )
  );

  defparam id01340.INIT = 16'h75AE;
  LUT4 id01340 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03838)
  );

  defparam id01341.INIT = 16'h7D00;
  LUT4 id01341 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03835),
    .O(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x0 )
  );

  defparam id01342.INIT = 16'h75AE;
  LUT4 id01342 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03835)
  );

  defparam id01343.INIT = 16'h00BE;
  LUT4 id01343 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03836),
    .O(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x0 )
  );

  defparam id01344.INIT = 16'hE817;
  LUT4 id01344 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03836)
  );

  defparam id01345.INIT = 16'h7D00;
  LUT4 id01345 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03825),
    .O(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x0 )
  );

  defparam id01346.INIT = 16'h75AE;
  LUT4 id01346 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03825)
  );

  defparam id01347.INIT = 16'h00BE;
  LUT4 id01347 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03826),
    .O(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x0 )
  );

  defparam id01348.INIT = 16'hE817;
  LUT4 id01348 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03826)
  );

  defparam id01349.INIT = 16'h00BE;
  LUT4 id01349 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03823),
    .O(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x0 )
  );

  defparam id01350.INIT = 16'hE817;
  LUT4 id01350 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03823)
  );

  defparam id01351.INIT = 16'h00BE;
  LUT4 id01351 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03824),
    .O(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x0 )
  );

  defparam id01352.INIT = 16'hE817;
  LUT4 id01352 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03824)
  );

  defparam id01353.INIT = 16'h7D00;
  LUT4 id01353 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03829),
    .O(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x0 )
  );

  defparam id01354.INIT = 16'h75AE;
  LUT4 id01354 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03829)
  );

  defparam id01355.INIT = 16'h7D00;
  LUT4 id01355 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03830),
    .O(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x0 )
  );

  defparam id01356.INIT = 16'h75AE;
  LUT4 id01356 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03830)
  );

  defparam id01357.INIT = 16'h7D00;
  LUT4 id01357 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03827),
    .O(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x0 )
  );

  defparam id01358.INIT = 16'h75AE;
  LUT4 id01358 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03827)
  );

  defparam id01359.INIT = 16'h7D00;
  LUT4 id01359 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03828),
    .O(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x0 )
  );

  defparam id01360.INIT = 16'h75AE;
  LUT4 id01360 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[24] ),
    .O(id03828)
  );

  defparam id01361.INIT = 16'h00BE;
  LUT4 id01361 (
    .ADR0(id03850),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03753),
    .O(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x0 )
  );

  defparam id01362.INIT = 16'hE817;
  LUT4 id01362 (
    .ADR0(\net_Buf-pad-multiplier[23] ),
    .ADR1(\net_Buf-pad-multiplier[24] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[25] ),
    .O(id03753)
  );

  defparam id01363.INIT = 16'hABD5;
  LUT4 id01363 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[23] ),
    .ADR2(\net_Buf-pad-multiplier[24] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x0 )
  );

  defparam id01364.INIT = 16'h1760;
  LUT4 id01364 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 )
  );

  defparam id01365.INIT = 16'h7D00;
  LUT4 id01365 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03751),
    .O(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 )
  );

  defparam id01366.INIT = 4'h6;
  LUT2 id01366 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .O(id03754)
  );

  defparam id01367.INIT = 16'h75AE;
  LUT4 id01367 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03751)
  );

  defparam id01368.INIT = 16'h7D00;
  LUT4 id01368 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03752),
    .O(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x1 )
  );

  defparam id01369.INIT = 16'h75AE;
  LUT4 id01369 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03752)
  );

  defparam id01370.INIT = 16'h7D00;
  LUT4 id01370 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03757),
    .O(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x1 )
  );

  defparam id01371.INIT = 16'h75AE;
  LUT4 id01371 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03757)
  );

  defparam id01372.INIT = 16'h7D00;
  LUT4 id01372 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03758),
    .O(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x1 )
  );

  defparam id01373.INIT = 16'h75AE;
  LUT4 id01373 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03758)
  );

  defparam id01374.INIT = 16'h7D00;
  LUT4 id01374 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03755),
    .O(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x1 )
  );

  defparam id01375.INIT = 16'h75AE;
  LUT4 id01375 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03755)
  );

  defparam id01376.INIT = 16'h7D00;
  LUT4 id01376 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03756),
    .O(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x1 )
  );

  defparam id01377.INIT = 16'h75AE;
  LUT4 id01377 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03756)
  );

  defparam id01378.INIT = 16'h7D00;
  LUT4 id01378 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03745),
    .O(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x1 )
  );

  defparam id01379.INIT = 16'h75AE;
  LUT4 id01379 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03745)
  );

  defparam id01380.INIT = 16'h7D00;
  LUT4 id01380 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03746),
    .O(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x1 )
  );

  defparam id01381.INIT = 16'h75AE;
  LUT4 id01381 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03746)
  );

  defparam id01382.INIT = 16'h7D00;
  LUT4 id01382 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03743),
    .O(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x1 )
  );

  defparam id01383.INIT = 16'h75AE;
  LUT4 id01383 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03743)
  );

  defparam id01384.INIT = 16'h7D00;
  LUT4 id01384 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03744),
    .O(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x1 )
  );

  defparam id01385.INIT = 16'h75AE;
  LUT4 id01385 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03744)
  );

  defparam id01386.INIT = 16'h7D00;
  LUT4 id01386 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03749),
    .O(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x1 )
  );

  defparam id01387.INIT = 16'h75AE;
  LUT4 id01387 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03749)
  );

  defparam id01388.INIT = 16'h7D00;
  LUT4 id01388 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03750),
    .O(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x1 )
  );

  defparam id01389.INIT = 16'h75AE;
  LUT4 id01389 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03750)
  );

  defparam id01390.INIT = 16'h00BE;
  LUT4 id01390 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03747),
    .O(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x1 )
  );

  defparam id01391.INIT = 16'hE817;
  LUT4 id01391 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(id03747)
  );

  defparam id01392.INIT = 16'h7D00;
  LUT4 id01392 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03748),
    .O(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x1 )
  );

  defparam id01393.INIT = 16'h75AE;
  LUT4 id01393 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03748)
  );

  defparam id01394.INIT = 16'h7D00;
  LUT4 id01394 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03737),
    .O(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x1 )
  );

  defparam id01395.INIT = 16'h75AE;
  LUT4 id01395 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03737)
  );

  defparam id01396.INIT = 16'h7D00;
  LUT4 id01396 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03738),
    .O(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x1 )
  );

  defparam id01397.INIT = 16'h75AE;
  LUT4 id01397 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03738)
  );

  defparam id01398.INIT = 16'h7D00;
  LUT4 id01398 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03735),
    .O(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x1 )
  );

  defparam id01399.INIT = 16'h75AE;
  LUT4 id01399 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03735)
  );

  defparam id01400.INIT = 16'h7D00;
  LUT4 id01400 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03736),
    .O(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x1 )
  );

  defparam id01401.INIT = 16'h75AE;
  LUT4 id01401 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03736)
  );

  defparam id01402.INIT = 16'h7D00;
  LUT4 id01402 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03741),
    .O(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x1 )
  );

  defparam id01403.INIT = 16'h75AE;
  LUT4 id01403 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03741)
  );

  defparam id01404.INIT = 16'h00BE;
  LUT4 id01404 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03742),
    .O(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x1 )
  );

  defparam id01405.INIT = 16'hE817;
  LUT4 id01405 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(id03742)
  );

  defparam id01406.INIT = 16'h7D00;
  LUT4 id01406 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03739),
    .O(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x1 )
  );

  defparam id01407.INIT = 16'h75AE;
  LUT4 id01407 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03739)
  );

  defparam id01408.INIT = 16'h7D00;
  LUT4 id01408 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03740),
    .O(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x1 )
  );

  defparam id01409.INIT = 16'h75AE;
  LUT4 id01409 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03740)
  );

  defparam id01410.INIT = 16'h7D00;
  LUT4 id01410 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03729),
    .O(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x1 )
  );

  defparam id01411.INIT = 16'h75AE;
  LUT4 id01411 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03729)
  );

  defparam id01412.INIT = 16'h7D00;
  LUT4 id01412 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03730),
    .O(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x1 )
  );

  defparam id01413.INIT = 16'h75AE;
  LUT4 id01413 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03730)
  );

  defparam id01414.INIT = 16'h7D00;
  LUT4 id01414 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03727),
    .O(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x1 )
  );

  defparam id01415.INIT = 16'h75AE;
  LUT4 id01415 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03727)
  );

  defparam id01416.INIT = 16'h7D00;
  LUT4 id01416 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03728),
    .O(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x1 )
  );

  defparam id01417.INIT = 16'h75AE;
  LUT4 id01417 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03728)
  );

  defparam id01418.INIT = 16'h7D00;
  LUT4 id01418 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03733),
    .O(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x1 )
  );

  defparam id01419.INIT = 16'h75AE;
  LUT4 id01419 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03733)
  );

  defparam id01420.INIT = 16'h00BE;
  LUT4 id01420 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03734),
    .O(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x1 )
  );

  defparam id01421.INIT = 16'hE817;
  LUT4 id01421 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(id03734)
  );

  defparam id01422.INIT = 16'h00BE;
  LUT4 id01422 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03731),
    .O(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x1 )
  );

  defparam id01423.INIT = 16'hE817;
  LUT4 id01423 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(id03731)
  );

  defparam id01424.INIT = 16'h7D00;
  LUT4 id01424 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03732),
    .O(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x1 )
  );

  defparam id01425.INIT = 16'h75AE;
  LUT4 id01425 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[26] ),
    .O(id03732)
  );

  defparam id01426.INIT = 16'h00BE;
  LUT4 id01426 (
    .ADR0(id03754),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03785),
    .O(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x1 )
  );

  defparam id01427.INIT = 16'hE817;
  LUT4 id01427 (
    .ADR0(\net_Buf-pad-multiplier[25] ),
    .ADR1(\net_Buf-pad-multiplier[26] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[27] ),
    .O(id03785)
  );

  defparam id01428.INIT = 16'hABD5;
  LUT4 id01428 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[25] ),
    .ADR2(\net_Buf-pad-multiplier[26] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x1 )
  );

  defparam id01429.INIT = 8'h78;
  LUT3 id01429 (
    .ADR0(\net_Buf-pad-multiplier[0] ),
    .ADR1(\net_Buf-pad-multiplicand[0] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .O(\u_compressor42_l0_0.CELLS[0].u_compressor42_cell.x0 )
  );

  defparam id01430.INIT = 16'h3C50;
  LUT4 id01430 (
    .ADR0(\net_Buf-pad-multiplicand[0] ),
    .ADR1(\net_Buf-pad-multiplicand[1] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 )
  );

  defparam id01431.INIT = 16'h3C50;
  LUT4 id01431 (
    .ADR0(\net_Buf-pad-multiplicand[1] ),
    .ADR1(\net_Buf-pad-multiplicand[2] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x0 )
  );

  defparam id01432.INIT = 16'h3C50;
  LUT4 id01432 (
    .ADR0(\net_Buf-pad-multiplicand[2] ),
    .ADR1(\net_Buf-pad-multiplicand[3] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x0 )
  );

  defparam id01433.INIT = 16'h3C50;
  LUT4 id01433 (
    .ADR0(\net_Buf-pad-multiplicand[3] ),
    .ADR1(\net_Buf-pad-multiplicand[4] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x0 )
  );

  defparam id01434.INIT = 16'h1760;
  LUT4 id01434 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x2 )
  );

  defparam id01435.INIT = 16'h00BE;
  LUT4 id01435 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id03783),
    .O(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x2 )
  );

  defparam id01436.INIT = 4'h6;
  LUT2 id01436 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .O(id03786)
  );

  defparam id01437.INIT = 16'hE817;
  LUT4 id01437 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03783)
  );

  defparam id01438.INIT = 16'h3C50;
  LUT4 id01438 (
    .ADR0(\net_Buf-pad-multiplicand[4] ),
    .ADR1(\net_Buf-pad-multiplicand[5] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x0 )
  );

  defparam id01439.INIT = 16'h00BE;
  LUT4 id01439 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03784),
    .O(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x2 )
  );

  defparam id01440.INIT = 16'hE817;
  LUT4 id01440 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03784)
  );

  defparam id01441.INIT = 16'h00BE;
  LUT4 id01441 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03789),
    .O(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x2 )
  );

  defparam id01442.INIT = 16'hE817;
  LUT4 id01442 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03789)
  );

  defparam id01443.INIT = 16'h00BE;
  LUT4 id01443 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03790),
    .O(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x2 )
  );

  defparam id01444.INIT = 16'hE817;
  LUT4 id01444 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03790)
  );

  defparam id01445.INIT = 16'h00BE;
  LUT4 id01445 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03787),
    .O(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x2 )
  );

  defparam id01446.INIT = 16'hE817;
  LUT4 id01446 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03787)
  );

  defparam id01447.INIT = 16'h00BE;
  LUT4 id01447 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03788),
    .O(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x2 )
  );

  defparam id01448.INIT = 16'hE817;
  LUT4 id01448 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03788)
  );

  defparam id01449.INIT = 16'h00BE;
  LUT4 id01449 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03777),
    .O(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x2 )
  );

  defparam id01450.INIT = 16'hE817;
  LUT4 id01450 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03777)
  );

  defparam id01451.INIT = 16'h00BE;
  LUT4 id01451 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03778),
    .O(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x2 )
  );

  defparam id01452.INIT = 16'hE817;
  LUT4 id01452 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03778)
  );

  defparam id01453.INIT = 16'h00BE;
  LUT4 id01453 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03775),
    .O(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x2 )
  );

  defparam id01454.INIT = 16'hE817;
  LUT4 id01454 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03775)
  );

  defparam id01455.INIT = 16'h00BE;
  LUT4 id01455 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03776),
    .O(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x2 )
  );

  defparam id01456.INIT = 16'hE817;
  LUT4 id01456 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03776)
  );

  defparam id01457.INIT = 16'h00BE;
  LUT4 id01457 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03781),
    .O(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x2 )
  );

  defparam id01458.INIT = 16'hE817;
  LUT4 id01458 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03781)
  );

  defparam id01459.INIT = 16'h3C50;
  LUT4 id01459 (
    .ADR0(\net_Buf-pad-multiplicand[5] ),
    .ADR1(\net_Buf-pad-multiplicand[6] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x0 )
  );

  defparam id01460.INIT = 16'h00BE;
  LUT4 id01460 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03782),
    .O(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x2 )
  );

  defparam id01461.INIT = 16'hE817;
  LUT4 id01461 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03782)
  );

  defparam id01462.INIT = 16'h00BE;
  LUT4 id01462 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03779),
    .O(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x2 )
  );

  defparam id01463.INIT = 16'hE817;
  LUT4 id01463 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03779)
  );

  defparam id01464.INIT = 16'h00BE;
  LUT4 id01464 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id03780),
    .O(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x2 )
  );

  defparam id01465.INIT = 16'hE817;
  LUT4 id01465 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03780)
  );

  defparam id01466.INIT = 16'h00BE;
  LUT4 id01466 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03769),
    .O(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x2 )
  );

  defparam id01467.INIT = 16'hE817;
  LUT4 id01467 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03769)
  );

  defparam id01468.INIT = 16'h00BE;
  LUT4 id01468 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03770),
    .O(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x2 )
  );

  defparam id01469.INIT = 16'hE817;
  LUT4 id01469 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03770)
  );

  defparam id01470.INIT = 16'h00BE;
  LUT4 id01470 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03767),
    .O(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x2 )
  );

  defparam id01471.INIT = 16'hE817;
  LUT4 id01471 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03767)
  );

  defparam id01472.INIT = 16'h00BE;
  LUT4 id01472 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03768),
    .O(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x2 )
  );

  defparam id01473.INIT = 16'hE817;
  LUT4 id01473 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03768)
  );

  defparam id01474.INIT = 16'h00BE;
  LUT4 id01474 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03773),
    .O(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x2 )
  );

  defparam id01475.INIT = 16'hE817;
  LUT4 id01475 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03773)
  );

  defparam id01476.INIT = 16'h00BE;
  LUT4 id01476 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03774),
    .O(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x2 )
  );

  defparam id01477.INIT = 16'hE817;
  LUT4 id01477 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03774)
  );

  defparam id01478.INIT = 16'h00BE;
  LUT4 id01478 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03771),
    .O(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x2 )
  );

  defparam id01479.INIT = 16'hE817;
  LUT4 id01479 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03771)
  );

  defparam id01480.INIT = 16'h3C50;
  LUT4 id01480 (
    .ADR0(\net_Buf-pad-multiplicand[6] ),
    .ADR1(\net_Buf-pad-multiplicand[7] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x0 )
  );

  defparam id01481.INIT = 16'h00BE;
  LUT4 id01481 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03772),
    .O(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x2 )
  );

  defparam id01482.INIT = 16'hE817;
  LUT4 id01482 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03772)
  );

  defparam id01483.INIT = 16'h00BE;
  LUT4 id01483 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03761),
    .O(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x2 )
  );

  defparam id01484.INIT = 16'hE817;
  LUT4 id01484 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03761)
  );

  defparam id01485.INIT = 16'h00BE;
  LUT4 id01485 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03762),
    .O(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x2 )
  );

  defparam id01486.INIT = 16'hE817;
  LUT4 id01486 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03762)
  );

  defparam id01487.INIT = 16'h00BE;
  LUT4 id01487 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03759),
    .O(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x2 )
  );

  defparam id01488.INIT = 16'hE817;
  LUT4 id01488 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03759)
  );

  defparam id01489.INIT = 16'h00BE;
  LUT4 id01489 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03760),
    .O(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x2 )
  );

  defparam id01490.INIT = 16'hE817;
  LUT4 id01490 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03760)
  );

  defparam id01491.INIT = 16'h00BE;
  LUT4 id01491 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03765),
    .O(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x2 )
  );

  defparam id01492.INIT = 16'hE817;
  LUT4 id01492 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03765)
  );

  defparam id01493.INIT = 16'h00BE;
  LUT4 id01493 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03766),
    .O(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x2 )
  );

  defparam id01494.INIT = 16'hE817;
  LUT4 id01494 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03766)
  );

  defparam id01495.INIT = 16'h00BE;
  LUT4 id01495 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03763),
    .O(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x2 )
  );

  defparam id01496.INIT = 16'hE817;
  LUT4 id01496 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03763)
  );

  defparam id01497.INIT = 16'h00BE;
  LUT4 id01497 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03764),
    .O(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x2 )
  );

  defparam id01498.INIT = 16'hE817;
  LUT4 id01498 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03764)
  );

  defparam id01499.INIT = 16'h00BE;
  LUT4 id01499 (
    .ADR0(id03786),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03945),
    .O(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x2 )
  );

  defparam id01500.INIT = 16'hE817;
  LUT4 id01500 (
    .ADR0(\net_Buf-pad-multiplier[27] ),
    .ADR1(\net_Buf-pad-multiplier[28] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[29] ),
    .O(id03945)
  );

  defparam id01501.INIT = 16'h3C50;
  LUT4 id01501 (
    .ADR0(\net_Buf-pad-multiplicand[7] ),
    .ADR1(\net_Buf-pad-multiplicand[8] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x0 )
  );

  defparam id01502.INIT = 16'hABD5;
  LUT4 id01502 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[27] ),
    .ADR2(\net_Buf-pad-multiplier[28] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x2 )
  );

  defparam id01503.INIT = 16'h3C50;
  LUT4 id01503 (
    .ADR0(\net_Buf-pad-multiplicand[8] ),
    .ADR1(\net_Buf-pad-multiplicand[9] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x0 )
  );

  defparam id01504.INIT = 16'h3C50;
  LUT4 id01504 (
    .ADR0(\net_Buf-pad-multiplicand[9] ),
    .ADR1(\net_Buf-pad-multiplicand[10] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x0 )
  );

  defparam id01505.INIT = 16'h3C50;
  LUT4 id01505 (
    .ADR0(\net_Buf-pad-multiplicand[10] ),
    .ADR1(\net_Buf-pad-multiplicand[11] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x0 )
  );

  defparam id01506.INIT = 16'h3C50;
  LUT4 id01506 (
    .ADR0(\net_Buf-pad-multiplicand[11] ),
    .ADR1(\net_Buf-pad-multiplicand[12] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x0 )
  );

  defparam id01507.INIT = 16'h3C50;
  LUT4 id01507 (
    .ADR0(\net_Buf-pad-multiplicand[12] ),
    .ADR1(\net_Buf-pad-multiplicand[13] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x0 )
  );

  defparam id01508.INIT = 16'h3C50;
  LUT4 id01508 (
    .ADR0(\net_Buf-pad-multiplicand[13] ),
    .ADR1(\net_Buf-pad-multiplicand[14] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x0 )
  );

  defparam id01509.INIT = 16'h3C50;
  LUT4 id01509 (
    .ADR0(\net_Buf-pad-multiplicand[14] ),
    .ADR1(\net_Buf-pad-multiplicand[15] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x0 )
  );

  defparam id01510.INIT = 16'h3C50;
  LUT4 id01510 (
    .ADR0(\net_Buf-pad-multiplicand[15] ),
    .ADR1(\net_Buf-pad-multiplicand[16] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x0 )
  );

  defparam id01511.INIT = 16'h3C50;
  LUT4 id01511 (
    .ADR0(\net_Buf-pad-multiplicand[16] ),
    .ADR1(\net_Buf-pad-multiplicand[17] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x0 )
  );

  defparam id01512.INIT = 16'h3C50;
  LUT4 id01512 (
    .ADR0(\net_Buf-pad-multiplicand[17] ),
    .ADR1(\net_Buf-pad-multiplicand[18] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x0 )
  );

  defparam id01513.INIT = 16'h3C50;
  LUT4 id01513 (
    .ADR0(\net_Buf-pad-multiplicand[18] ),
    .ADR1(\net_Buf-pad-multiplicand[19] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x0 )
  );

  defparam id01514.INIT = 16'h3C50;
  LUT4 id01514 (
    .ADR0(\net_Buf-pad-multiplicand[19] ),
    .ADR1(\net_Buf-pad-multiplicand[20] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x0 )
  );

  defparam id01515.INIT = 16'h3C50;
  LUT4 id01515 (
    .ADR0(\net_Buf-pad-multiplicand[20] ),
    .ADR1(\net_Buf-pad-multiplicand[21] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x0 )
  );

  defparam id01516.INIT = 16'h3C50;
  LUT4 id01516 (
    .ADR0(\net_Buf-pad-multiplicand[21] ),
    .ADR1(\net_Buf-pad-multiplicand[22] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x0 )
  );

  defparam id01517.INIT = 16'h3C50;
  LUT4 id01517 (
    .ADR0(\net_Buf-pad-multiplicand[22] ),
    .ADR1(\net_Buf-pad-multiplicand[23] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x0 )
  );

  defparam id01518.INIT = 16'h3C50;
  LUT4 id01518 (
    .ADR0(\net_Buf-pad-multiplicand[23] ),
    .ADR1(\net_Buf-pad-multiplicand[24] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x0 )
  );

  defparam id01519.INIT = 16'h3C50;
  LUT4 id01519 (
    .ADR0(\net_Buf-pad-multiplicand[24] ),
    .ADR1(\net_Buf-pad-multiplicand[25] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x0 )
  );

  defparam id01520.INIT = 16'h3C50;
  LUT4 id01520 (
    .ADR0(\net_Buf-pad-multiplicand[25] ),
    .ADR1(\net_Buf-pad-multiplicand[26] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x0 )
  );

  defparam id01521.INIT = 16'h1760;
  LUT4 id01521 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x3 )
  );

  defparam id01522.INIT = 16'hBEAA;
  LUT4 id01522 (
    .ADR0(id03946),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x3 )
  );

  defparam id01523.INIT = 4'h6;
  LUT2 id01523 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .O(id03944)
  );

  defparam id01524.INIT = 8'h70;
  LUT3 id01524 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplier[29] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03943)
  );

  defparam id01525.INIT = 16'h0180;
  LUT4 id01525 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03946)
  );

  defparam id01526.INIT = 16'h3CAA;
  LUT4 id01526 (
    .ADR0(id03949),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x3 )
  );

  defparam id01527.INIT = 8'h18;
  LUT3 id01527 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[1] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03949)
  );

  defparam id01528.INIT = 16'h3C50;
  LUT4 id01528 (
    .ADR0(\net_Buf-pad-multiplicand[26] ),
    .ADR1(\net_Buf-pad-multiplicand[27] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x0 )
  );

  defparam id01529.INIT = 16'h3CAA;
  LUT4 id01529 (
    .ADR0(id03950),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[11].u_compressor42_cell.x3 )
  );

  defparam id01530.INIT = 8'h18;
  LUT3 id01530 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[2] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03950)
  );

  defparam id01531.INIT = 16'h3CAA;
  LUT4 id01531 (
    .ADR0(id03947),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[12].u_compressor42_cell.x3 )
  );

  defparam id01532.INIT = 8'h18;
  LUT3 id01532 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[3] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03947)
  );

  defparam id01533.INIT = 16'h3CAA;
  LUT4 id01533 (
    .ADR0(id03948),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[13].u_compressor42_cell.x3 )
  );

  defparam id01534.INIT = 8'h18;
  LUT3 id01534 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[4] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03948)
  );

  defparam id01535.INIT = 16'h3CAA;
  LUT4 id01535 (
    .ADR0(id03937),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[14].u_compressor42_cell.x3 )
  );

  defparam id01536.INIT = 8'h18;
  LUT3 id01536 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[5] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03937)
  );

  defparam id01537.INIT = 16'h3CAA;
  LUT4 id01537 (
    .ADR0(id03938),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[15].u_compressor42_cell.x3 )
  );

  defparam id01538.INIT = 8'h18;
  LUT3 id01538 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[6] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03938)
  );

  defparam id01539.INIT = 16'h3CAA;
  LUT4 id01539 (
    .ADR0(id03935),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[16].u_compressor42_cell.x3 )
  );

  defparam id01540.INIT = 8'h18;
  LUT3 id01540 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[7] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03935)
  );

  defparam id01541.INIT = 16'h3CAA;
  LUT4 id01541 (
    .ADR0(id03936),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[17].u_compressor42_cell.x3 )
  );

  defparam id01542.INIT = 8'h18;
  LUT3 id01542 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[8] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03936)
  );

  defparam id01543.INIT = 16'h3CAA;
  LUT4 id01543 (
    .ADR0(id03941),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[18].u_compressor42_cell.x3 )
  );

  defparam id01544.INIT = 8'h18;
  LUT3 id01544 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[9] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03941)
  );

  defparam id01545.INIT = 16'h3CAA;
  LUT4 id01545 (
    .ADR0(id03942),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[19].u_compressor42_cell.x3 )
  );

  defparam id01546.INIT = 8'h18;
  LUT3 id01546 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[10] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03942)
  );

  defparam id01547.INIT = 16'h3CAA;
  LUT4 id01547 (
    .ADR0(id03939),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[20].u_compressor42_cell.x3 )
  );

  defparam id01548.INIT = 8'h18;
  LUT3 id01548 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[11] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03939)
  );

  defparam id01549.INIT = 16'h3C50;
  LUT4 id01549 (
    .ADR0(\net_Buf-pad-multiplicand[27] ),
    .ADR1(\net_Buf-pad-multiplicand[28] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x0 )
  );

  defparam id01550.INIT = 16'h3CAA;
  LUT4 id01550 (
    .ADR0(id03940),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[21].u_compressor42_cell.x3 )
  );

  defparam id01551.INIT = 8'h18;
  LUT3 id01551 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[12] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03940)
  );

  defparam id01552.INIT = 16'h3CAA;
  LUT4 id01552 (
    .ADR0(id03929),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[22].u_compressor42_cell.x3 )
  );

  defparam id01553.INIT = 8'h18;
  LUT3 id01553 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[13] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03929)
  );

  defparam id01554.INIT = 16'h3CAA;
  LUT4 id01554 (
    .ADR0(id03930),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[23].u_compressor42_cell.x3 )
  );

  defparam id01555.INIT = 8'h18;
  LUT3 id01555 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[14] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03930)
  );

  defparam id01556.INIT = 16'h3CAA;
  LUT4 id01556 (
    .ADR0(id03927),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[24].u_compressor42_cell.x3 )
  );

  defparam id01557.INIT = 8'h18;
  LUT3 id01557 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[15] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03927)
  );

  defparam id01558.INIT = 16'h3CAA;
  LUT4 id01558 (
    .ADR0(id03928),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[25].u_compressor42_cell.x3 )
  );

  defparam id01559.INIT = 8'h18;
  LUT3 id01559 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[16] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03928)
  );

  defparam id01560.INIT = 16'h3CAA;
  LUT4 id01560 (
    .ADR0(id03933),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03944),
    .O(\u_compressor42_l0_3.CELLS[26].u_compressor42_cell.x3 )
  );

  defparam id01561.INIT = 8'h18;
  LUT3 id01561 (
    .ADR0(\net_Buf-pad-multiplier[30] ),
    .ADR1(\net_Buf-pad-multiplicand[17] ),
    .ADR2(\net_Buf-pad-multiplier[31] ),
    .O(id03933)
  );

  defparam id01562.INIT = 16'h00BE;
  LUT4 id01562 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03934),
    .O(\u_compressor42_l0_3.CELLS[27].u_compressor42_cell.x3 )
  );

  defparam id01563.INIT = 16'hE817;
  LUT4 id01563 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03934)
  );

  defparam id01564.INIT = 16'h00BE;
  LUT4 id01564 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03931),
    .O(\u_compressor42_l0_3.CELLS[28].u_compressor42_cell.x3 )
  );

  defparam id01565.INIT = 16'hE817;
  LUT4 id01565 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03931)
  );

  defparam id01566.INIT = 16'h00BE;
  LUT4 id01566 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03932),
    .O(\u_compressor42_l0_3.CELLS[29].u_compressor42_cell.x3 )
  );

  defparam id01567.INIT = 16'hE817;
  LUT4 id01567 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03932)
  );

  defparam id01568.INIT = 16'h00BE;
  LUT4 id01568 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03921),
    .O(\u_compressor42_l0_3.CELLS[30].u_compressor42_cell.x3 )
  );

  defparam id01569.INIT = 16'hE817;
  LUT4 id01569 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03921)
  );

  defparam id01570.INIT = 16'h3C50;
  LUT4 id01570 (
    .ADR0(\net_Buf-pad-multiplicand[28] ),
    .ADR1(\net_Buf-pad-multiplicand[29] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x0 )
  );

  defparam id01571.INIT = 16'h00BE;
  LUT4 id01571 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03922),
    .O(\u_compressor42_l0_3.CELLS[31].u_compressor42_cell.x3 )
  );

  defparam id01572.INIT = 16'hE817;
  LUT4 id01572 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03922)
  );

  defparam id01573.INIT = 16'h00BE;
  LUT4 id01573 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03919),
    .O(\u_compressor42_l0_3.CELLS[32].u_compressor42_cell.x3 )
  );

  defparam id01574.INIT = 16'hE817;
  LUT4 id01574 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03919)
  );

  defparam id01575.INIT = 16'h00BE;
  LUT4 id01575 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03920),
    .O(\u_compressor42_l0_3.CELLS[33].u_compressor42_cell.x3 )
  );

  defparam id01576.INIT = 16'hE817;
  LUT4 id01576 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03920)
  );

  defparam id01577.INIT = 16'h00BE;
  LUT4 id01577 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03925),
    .O(\u_compressor42_l0_3.CELLS[34].u_compressor42_cell.x3 )
  );

  defparam id01578.INIT = 16'hE817;
  LUT4 id01578 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03925)
  );

  defparam id01579.INIT = 16'h00BE;
  LUT4 id01579 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03926),
    .O(\u_compressor42_l0_3.CELLS[35].u_compressor42_cell.x3 )
  );

  defparam id01580.INIT = 16'hE817;
  LUT4 id01580 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03926)
  );

  defparam id01581.INIT = 16'h00BE;
  LUT4 id01581 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03923),
    .O(\u_compressor42_l0_3.CELLS[36].u_compressor42_cell.x3 )
  );

  defparam id01582.INIT = 16'hE817;
  LUT4 id01582 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03923)
  );

  defparam id01583.INIT = 16'h00BE;
  LUT4 id01583 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03924),
    .O(\u_compressor42_l0_3.CELLS[37].u_compressor42_cell.x3 )
  );

  defparam id01584.INIT = 16'hE817;
  LUT4 id01584 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03924)
  );

  defparam id01585.INIT = 16'h00BE;
  LUT4 id01585 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03977),
    .O(\u_compressor42_l0_3.CELLS[38].u_compressor42_cell.x3 )
  );

  defparam id01586.INIT = 16'hE817;
  LUT4 id01586 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03977)
  );

  defparam id01587.INIT = 16'h00BE;
  LUT4 id01587 (
    .ADR0(id03944),
    .ADR1(id03943),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03978),
    .O(\u_compressor42_l0_3.CELLS[39].u_compressor42_cell.x3 )
  );

  defparam id01588.INIT = 16'hE817;
  LUT4 id01588 (
    .ADR0(\net_Buf-pad-multiplier[29] ),
    .ADR1(\net_Buf-pad-multiplier[30] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[31] ),
    .O(id03978)
  );

  defparam id01589.INIT = 16'hABD5;
  LUT4 id01589 (
    .ADR0(\net_Buf-pad-multiplier[31] ),
    .ADR1(\net_Buf-pad-multiplier[29] ),
    .ADR2(\net_Buf-pad-multiplier[30] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_3.CELLS[40].u_compressor42_cell.x3 )
  );

  defparam id01590.INIT = 16'h3C50;
  LUT4 id01590 (
    .ADR0(\net_Buf-pad-multiplicand[29] ),
    .ADR1(\net_Buf-pad-multiplicand[30] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x0 )
  );

  defparam id01591.INIT = 16'h3C50;
  LUT4 id01591 (
    .ADR0(\net_Buf-pad-multiplicand[30] ),
    .ADR1(\net_Buf-pad-multiplicand[31] ),
    .ADR2(\net_Buf-pad-multiplier[1] ),
    .ADR3(\net_Buf-pad-multiplier[0] ),
    .O(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x0 )
  );

  defparam id01592.INIT = 8'h2C;
  LUT3 id01592 (
    .ADR0(\net_Buf-pad-multiplier[0] ),
    .ADR1(\net_Buf-pad-multiplier[1] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x0 )
  );

  defparam id01593.INIT = 16'h1760;
  LUT4 id01593 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x1 )
  );

  defparam id01594.INIT = 16'h00BE;
  LUT4 id01594 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(id03976),
    .O(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 )
  );

  defparam id01595.INIT = 4'h6;
  LUT2 id01595 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .O(id03975)
  );

  defparam id01596.INIT = 16'hE817;
  LUT4 id01596 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03976)
  );

  defparam id01597.INIT = 16'h00BE;
  LUT4 id01597 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03981),
    .O(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x1 )
  );

  defparam id01598.INIT = 16'hE817;
  LUT4 id01598 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03981)
  );

  defparam id01599.INIT = 16'h00BE;
  LUT4 id01599 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03982),
    .O(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x1 )
  );

  defparam id01600.INIT = 16'hE817;
  LUT4 id01600 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03982)
  );

  defparam id01601.INIT = 16'h00BE;
  LUT4 id01601 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(id03979),
    .O(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x1 )
  );

  defparam id01602.INIT = 16'hE817;
  LUT4 id01602 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03979)
  );

  defparam id01603.INIT = 16'h00BE;
  LUT4 id01603 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03980),
    .O(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x1 )
  );

  defparam id01604.INIT = 16'hE817;
  LUT4 id01604 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03980)
  );

  defparam id01605.INIT = 16'h00BE;
  LUT4 id01605 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03969),
    .O(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x1 )
  );

  defparam id01606.INIT = 16'hE817;
  LUT4 id01606 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03969)
  );

  defparam id01607.INIT = 16'h00BE;
  LUT4 id01607 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03970),
    .O(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x1 )
  );

  defparam id01608.INIT = 16'hE817;
  LUT4 id01608 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03970)
  );

  defparam id01609.INIT = 16'h00BE;
  LUT4 id01609 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(id03967),
    .O(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x1 )
  );

  defparam id01610.INIT = 16'hE817;
  LUT4 id01610 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03967)
  );

  defparam id01611.INIT = 16'h00BE;
  LUT4 id01611 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03968),
    .O(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x1 )
  );

  defparam id01612.INIT = 16'hE817;
  LUT4 id01612 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03968)
  );

  defparam id01613.INIT = 16'h00BE;
  LUT4 id01613 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03973),
    .O(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x1 )
  );

  defparam id01614.INIT = 16'hE817;
  LUT4 id01614 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03973)
  );

  defparam id01615.INIT = 16'h00BE;
  LUT4 id01615 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03974),
    .O(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x1 )
  );

  defparam id01616.INIT = 16'hE817;
  LUT4 id01616 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03974)
  );

  defparam id01617.INIT = 16'h00BE;
  LUT4 id01617 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03971),
    .O(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x1 )
  );

  defparam id01618.INIT = 16'hE817;
  LUT4 id01618 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03971)
  );

  defparam id01619.INIT = 16'h00BE;
  LUT4 id01619 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(id03972),
    .O(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x1 )
  );

  defparam id01620.INIT = 16'hE817;
  LUT4 id01620 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03972)
  );

  defparam id01621.INIT = 16'h00BE;
  LUT4 id01621 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id03961),
    .O(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x1 )
  );

  defparam id01622.INIT = 16'hE817;
  LUT4 id01622 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03961)
  );

  defparam id01623.INIT = 16'h00BE;
  LUT4 id01623 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03962),
    .O(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x1 )
  );

  defparam id01624.INIT = 16'hE817;
  LUT4 id01624 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03962)
  );

  defparam id01625.INIT = 16'h00BE;
  LUT4 id01625 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03959),
    .O(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x1 )
  );

  defparam id01626.INIT = 16'hE817;
  LUT4 id01626 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03959)
  );

  defparam id01627.INIT = 16'h00BE;
  LUT4 id01627 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(id03960),
    .O(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x1 )
  );

  defparam id01628.INIT = 16'hE817;
  LUT4 id01628 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03960)
  );

  defparam id01629.INIT = 16'h00BE;
  LUT4 id01629 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03965),
    .O(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x1 )
  );

  defparam id01630.INIT = 16'hE817;
  LUT4 id01630 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03965)
  );

  defparam id01631.INIT = 16'h00BE;
  LUT4 id01631 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03966),
    .O(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x1 )
  );

  defparam id01632.INIT = 16'hE817;
  LUT4 id01632 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03966)
  );

  defparam id01633.INIT = 16'h00BE;
  LUT4 id01633 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03963),
    .O(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x1 )
  );

  defparam id01634.INIT = 16'hE817;
  LUT4 id01634 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03963)
  );

  defparam id01635.INIT = 16'h00BE;
  LUT4 id01635 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03964),
    .O(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x1 )
  );

  defparam id01636.INIT = 16'hE817;
  LUT4 id01636 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03964)
  );

  defparam id01637.INIT = 16'h00BE;
  LUT4 id01637 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03953),
    .O(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x1 )
  );

  defparam id01638.INIT = 16'hE817;
  LUT4 id01638 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03953)
  );

  defparam id01639.INIT = 16'h00BE;
  LUT4 id01639 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03954),
    .O(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x1 )
  );

  defparam id01640.INIT = 16'hE817;
  LUT4 id01640 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03954)
  );

  defparam id01641.INIT = 16'h00BE;
  LUT4 id01641 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03951),
    .O(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x1 )
  );

  defparam id01642.INIT = 16'hE817;
  LUT4 id01642 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03951)
  );

  defparam id01643.INIT = 16'h00BE;
  LUT4 id01643 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03952),
    .O(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x1 )
  );

  defparam id01644.INIT = 16'hE817;
  LUT4 id01644 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03952)
  );

  defparam id01645.INIT = 16'h00BE;
  LUT4 id01645 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(id03957),
    .O(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x1 )
  );

  defparam id01646.INIT = 16'hE817;
  LUT4 id01646 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03957)
  );

  defparam id01647.INIT = 16'h00BE;
  LUT4 id01647 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03958),
    .O(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x1 )
  );

  defparam id01648.INIT = 16'hE817;
  LUT4 id01648 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03958)
  );

  defparam id01649.INIT = 16'h00BE;
  LUT4 id01649 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03955),
    .O(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x1 )
  );

  defparam id01650.INIT = 16'hE817;
  LUT4 id01650 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03955)
  );

  defparam id01651.INIT = 16'h00BE;
  LUT4 id01651 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03956),
    .O(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x1 )
  );

  defparam id01652.INIT = 16'hE817;
  LUT4 id01652 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03956)
  );

  defparam id01653.INIT = 16'h00BE;
  LUT4 id01653 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03881),
    .O(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x1 )
  );

  defparam id01654.INIT = 16'hE817;
  LUT4 id01654 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03881)
  );

  defparam id01655.INIT = 16'h00BE;
  LUT4 id01655 (
    .ADR0(id03975),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03882),
    .O(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x1 )
  );

  defparam id01656.INIT = 16'hE817;
  LUT4 id01656 (
    .ADR0(\net_Buf-pad-multiplier[1] ),
    .ADR1(\net_Buf-pad-multiplier[2] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[3] ),
    .O(id03882)
  );

  defparam id01657.INIT = 16'hABD5;
  LUT4 id01657 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[1] ),
    .ADR2(\net_Buf-pad-multiplier[2] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x1 )
  );

  defparam id01658.INIT = 16'h1760;
  LUT4 id01658 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x2 )
  );

  defparam id01659.INIT = 16'h7D00;
  LUT4 id01659 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(id03880),
    .O(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x2 )
  );

  defparam id01660.INIT = 4'h6;
  LUT2 id01660 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .O(id03879)
  );

  defparam id01661.INIT = 16'h75AE;
  LUT4 id01661 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03880)
  );

  defparam id01662.INIT = 16'h7D00;
  LUT4 id01662 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03885),
    .O(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x2 )
  );

  defparam id01663.INIT = 16'h75AE;
  LUT4 id01663 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[1] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03885)
  );

  defparam id01664.INIT = 16'h00BE;
  LUT4 id01664 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[2] ),
    .ADR3(id03886),
    .O(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x2 )
  );

  defparam id01665.INIT = 16'hE817;
  LUT4 id01665 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03886)
  );

  defparam id01666.INIT = 16'h7D00;
  LUT4 id01666 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03883),
    .O(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x2 )
  );

  defparam id01667.INIT = 16'h75AE;
  LUT4 id01667 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[3] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03883)
  );

  defparam id01668.INIT = 16'h00BE;
  LUT4 id01668 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[4] ),
    .ADR3(id03884),
    .O(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x2 )
  );

  defparam id01669.INIT = 16'hE817;
  LUT4 id01669 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03884)
  );

  defparam id01670.INIT = 16'h00BE;
  LUT4 id01670 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[5] ),
    .ADR3(id03873),
    .O(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x2 )
  );

  defparam id01671.INIT = 16'hE817;
  LUT4 id01671 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03873)
  );

  defparam id01672.INIT = 16'h00BE;
  LUT4 id01672 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[6] ),
    .ADR3(id03874),
    .O(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x2 )
  );

  defparam id01673.INIT = 16'hE817;
  LUT4 id01673 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03874)
  );

  defparam id01674.INIT = 16'h7D00;
  LUT4 id01674 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(id03871),
    .O(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x2 )
  );

  defparam id01675.INIT = 16'h75AE;
  LUT4 id01675 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[7] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03871)
  );

  defparam id01676.INIT = 16'h7D00;
  LUT4 id01676 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(id03872),
    .O(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x2 )
  );

  defparam id01677.INIT = 16'h75AE;
  LUT4 id01677 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[8] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03872)
  );

  defparam id01678.INIT = 16'h7D00;
  LUT4 id01678 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(id03877),
    .O(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x2 )
  );

  defparam id01679.INIT = 16'h75AE;
  LUT4 id01679 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[9] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03877)
  );

  defparam id01680.INIT = 16'h7D00;
  LUT4 id01680 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03878),
    .O(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x2 )
  );

  defparam id01681.INIT = 16'h75AE;
  LUT4 id01681 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[10] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03878)
  );

  defparam id01682.INIT = 16'h00BE;
  LUT4 id01682 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[11] ),
    .ADR3(id03875),
    .O(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x2 )
  );

  defparam id01683.INIT = 16'hE817;
  LUT4 id01683 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03875)
  );

  defparam id01684.INIT = 16'h7D00;
  LUT4 id01684 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(id03876),
    .O(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x2 )
  );

  defparam id01685.INIT = 16'h75AE;
  LUT4 id01685 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[12] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03876)
  );

  defparam id01686.INIT = 16'h7D00;
  LUT4 id01686 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(id03865),
    .O(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x2 )
  );

  defparam id01687.INIT = 16'h75AE;
  LUT4 id01687 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[13] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03865)
  );

  defparam id01688.INIT = 16'h7D00;
  LUT4 id01688 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03866),
    .O(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x2 )
  );

  defparam id01689.INIT = 16'h75AE;
  LUT4 id01689 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[14] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03866)
  );

  defparam id01690.INIT = 16'h00BE;
  LUT4 id01690 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[15] ),
    .ADR3(id03863),
    .O(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x2 )
  );

  defparam id01691.INIT = 16'hE817;
  LUT4 id01691 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03863)
  );

  defparam id01692.INIT = 16'h7D00;
  LUT4 id01692 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(id03864),
    .O(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x2 )
  );

  defparam id01693.INIT = 16'h75AE;
  LUT4 id01693 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[16] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03864)
  );

  defparam id01694.INIT = 16'h7D00;
  LUT4 id01694 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(id03869),
    .O(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x2 )
  );

  defparam id01695.INIT = 16'h75AE;
  LUT4 id01695 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[17] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03869)
  );

  defparam id01696.INIT = 16'h7D00;
  LUT4 id01696 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(id03870),
    .O(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x2 )
  );

  defparam id01697.INIT = 16'h75AE;
  LUT4 id01697 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[18] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03870)
  );

  defparam id01698.INIT = 16'h7D00;
  LUT4 id01698 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(id03867),
    .O(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x2 )
  );

  defparam id01699.INIT = 16'h75AE;
  LUT4 id01699 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[19] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03867)
  );

  defparam id01700.INIT = 16'h7D00;
  LUT4 id01700 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(id03868),
    .O(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x2 )
  );

  defparam id01701.INIT = 16'h75AE;
  LUT4 id01701 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[20] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03868)
  );

  defparam id01702.INIT = 16'h7D00;
  LUT4 id01702 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(id03857),
    .O(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x2 )
  );

  defparam id01703.INIT = 16'h75AE;
  LUT4 id01703 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[21] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03857)
  );

  defparam id01704.INIT = 16'h7D00;
  LUT4 id01704 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(id03858),
    .O(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x2 )
  );

  defparam id01705.INIT = 16'h75AE;
  LUT4 id01705 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[22] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03858)
  );

  defparam id01706.INIT = 16'h7D00;
  LUT4 id01706 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03855),
    .O(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x2 )
  );

  defparam id01707.INIT = 16'h75AE;
  LUT4 id01707 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[23] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03855)
  );

  defparam id01708.INIT = 16'h00BE;
  LUT4 id01708 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[24] ),
    .ADR3(id03856),
    .O(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x2 )
  );

  defparam id01709.INIT = 16'hE817;
  LUT4 id01709 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03856)
  );

  defparam id01710.INIT = 16'h7D00;
  LUT4 id01710 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(id03861),
    .O(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x2 )
  );

  defparam id01711.INIT = 16'h75AE;
  LUT4 id01711 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[25] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03861)
  );

  defparam id01712.INIT = 16'h7D00;
  LUT4 id01712 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03862),
    .O(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x2 )
  );

  defparam id01713.INIT = 16'h75AE;
  LUT4 id01713 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[5] ),
    .ADR2(\net_Buf-pad-multiplicand[26] ),
    .ADR3(\net_Buf-pad-multiplier[4] ),
    .O(id03862)
  );

  defparam id01714.INIT = 16'h00BE;
  LUT4 id01714 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[27] ),
    .ADR3(id03859),
    .O(\u_compressor42_l0_0.CELLS[32].u_compressor42_cell.x2 )
  );

  defparam id01715.INIT = 16'hE817;
  LUT4 id01715 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03859)
  );

  defparam id01716.INIT = 16'h00BE;
  LUT4 id01716 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[28] ),
    .ADR3(id03860),
    .O(\u_compressor42_l0_0.CELLS[33].u_compressor42_cell.x2 )
  );

  defparam id01717.INIT = 16'hE817;
  LUT4 id01717 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03860)
  );

  defparam id01718.INIT = 16'h00BE;
  LUT4 id01718 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[29] ),
    .ADR3(id03913),
    .O(\u_compressor42_l0_0.CELLS[34].u_compressor42_cell.x2 )
  );

  defparam id01719.INIT = 16'hE817;
  LUT4 id01719 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03913)
  );

  defparam id01720.INIT = 16'h00BE;
  LUT4 id01720 (
    .ADR0(id03879),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\net_Buf-pad-multiplicand[30] ),
    .ADR3(id03914),
    .O(\u_compressor42_l0_0.CELLS[35].u_compressor42_cell.x2 )
  );

  defparam id01721.INIT = 16'hE817;
  LUT4 id01721 (
    .ADR0(\net_Buf-pad-multiplier[3] ),
    .ADR1(\net_Buf-pad-multiplier[4] ),
    .ADR2(\net_Buf-pad-multiplicand[31] ),
    .ADR3(\net_Buf-pad-multiplier[5] ),
    .O(id03914)
  );

  defparam id01722.INIT = 16'hABD5;
  LUT4 id01722 (
    .ADR0(\net_Buf-pad-multiplier[5] ),
    .ADR1(\net_Buf-pad-multiplier[3] ),
    .ADR2(\net_Buf-pad-multiplier[4] ),
    .ADR3(\net_Buf-pad-multiplicand[31] ),
    .O(\u_compressor42_l0_0.CELLS[36].u_compressor42_cell.x2 )
  );

  defparam id01723.INIT = 16'h1760;
  LUT4 id01723 (
    .ADR0(\net_Buf-pad-multiplier[5] ),
    .ADR1(\net_Buf-pad-multiplier[6] ),
    .ADR2(\net_Buf-pad-multiplicand[0] ),
    .ADR3(\net_Buf-pad-multiplier[7] ),
    .O(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x3 )
  );

  defparam id01724.INIT = 4'h1;
  LUT2 id01724 (
    .ADR0(id03911),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x3 )
  );

  defparam id01725.INIT = 16'hAC53;
  LUT4 id01725 (
    .ADR0(\net_Buf-pad-multiplicand[1] ),
    .ADR1(\net_Buf-pad-multiplicand[0] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03911)
  );

  defparam id01726.INIT = 4'h1;
  LUT2 id01726 (
    .ADR0(id03912),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x3 )
  );

  defparam id01727.INIT = 16'hAC53;
  LUT4 id01727 (
    .ADR0(\net_Buf-pad-multiplicand[2] ),
    .ADR1(\net_Buf-pad-multiplicand[1] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03912)
  );

  defparam id01728.INIT = 4'h1;
  LUT2 id01728 (
    .ADR0(id03917),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x3 )
  );

  defparam id01729.INIT = 16'hAC53;
  LUT4 id01729 (
    .ADR0(\net_Buf-pad-multiplicand[3] ),
    .ADR1(\net_Buf-pad-multiplicand[2] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03917)
  );

  defparam id01730.INIT = 4'h1;
  LUT2 id01730 (
    .ADR0(id03918),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x3 )
  );

  defparam id01731.INIT = 16'hAC53;
  LUT4 id01731 (
    .ADR0(\net_Buf-pad-multiplicand[4] ),
    .ADR1(\net_Buf-pad-multiplicand[3] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03918)
  );

  defparam id01732.INIT = 4'h1;
  LUT2 id01732 (
    .ADR0(id03915),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x3 )
  );

  defparam id01733.INIT = 16'hAC53;
  LUT4 id01733 (
    .ADR0(\net_Buf-pad-multiplicand[5] ),
    .ADR1(\net_Buf-pad-multiplicand[4] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03915)
  );

  defparam id01734.INIT = 4'h1;
  LUT2 id01734 (
    .ADR0(id03916),
    .ADR1(id04321),
    .O(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x3 )
  );

  defparam id01735.INIT = 16'hAC53;
  LUT4 id01735 (
    .ADR0(\net_Buf-pad-multiplicand[6] ),
    .ADR1(\net_Buf-pad-multiplicand[5] ),
    .ADR2(id04322),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id03916)
  );

  defparam id01736.INIT = 4'h6;
  LUT2 id01736 (
    .ADR0(\u_compressor42_l0_0.CELLS[0].u_compressor42_cell.x0 ),
    .ADR1(\net_Buf-pad-multiplier[1] ),
    .O(\net_Buf-pad-result[0] )
  );

  defparam id01737.INIT = 16'h8778;
  LUT4 id01737 (
    .ADR0(\u_compressor42_l0_0.CELLS[0].u_compressor42_cell.x0 ),
    .ADR1(\net_Buf-pad-multiplier[1] ),
    .ADR2(\u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(\net_Buf-pad-result[1] )
  );

  defparam id01738.INIT = 16'h07F8;
  LUT4 id01738 (
    .ADR0(\u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(id03905),
    .ADR3(id03906),
    .O(\net_Buf-pad-result[2] )
  );

  defparam id01739.INIT = 16'h6000;
  LUT4 id01739 (
    .ADR0(\u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[0].u_compressor42_cell.x0 ),
    .ADR3(\net_Buf-pad-multiplier[1] ),
    .O(id03905)
  );

  defparam id01740.INIT = 8'h96;
  LUT3 id01740 (
    .ADR0(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x1 ),
    .O(id03906)
  );

  defparam id01741.INIT = 16'h9669;
  LUT4 id01741 (
    .ADR0(id03903),
    .ADR1(id03904),
    .ADR2(id03909),
    .ADR3(id03910),
    .O(\net_Buf-pad-result[3] )
  );

  defparam id01742.INIT = 8'h80;
  LUT3 id01742 (
    .ADR0(id03906),
    .ADR1(\u_compressor42_l0_0.CELLS[1].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .O(id03903)
  );

  defparam id01743.INIT = 4'h8;
  LUT2 id01743 (
    .ADR0(id03905),
    .ADR1(id03906),
    .O(id03904)
  );

  defparam id01744.INIT = 4'h1;
  LUT2 id01744 (
    .ADR0(id03907),
    .ADR1(id03908),
    .O(id03909)
  );

  defparam id01745.INIT = 4'h8;
  LUT2 id01745 (
    .ADR0(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x1 ),
    .O(id03907)
  );

  defparam id01746.INIT = 8'h60;
  LUT3 id01746 (
    .ADR0(\DECODE_GEN[1].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[2].u_compressor42_cell.x0 ),
    .O(id03908)
  );

  defparam id01747.INIT = 8'h96;
  LUT3 id01747 (
    .ADR0(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ),
    .O(id03910)
  );

  defparam id01748.INIT = 4'h9;
  LUT2 id01748 (
    .ADR0(id03897),
    .ADR1(id03898),
    .O(\net_Buf-pad-result[5] )
  );

  defparam id01749.INIT = 16'h32F3;
  LUT4 id01749 (
    .ADR0(id03908),
    .ADR1(id03895),
    .ADR2(id03896),
    .ADR3(id03901),
    .O(id03897)
  );

  defparam id01750.INIT = 8'h90;
  LUT3 id01750 (
    .ADR0(id03909),
    .ADR1(id03910),
    .ADR2(id03904),
    .O(id03895)
  );

  defparam id01751.INIT = 16'h7887;
  LUT4 id01751 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ),
    .ADR2(id03902),
    .ADR3(id03899),
    .O(id03901)
  );

  defparam id01752.INIT = 16'h8EE8;
  LUT4 id01752 (
    .ADR0(id03907),
    .ADR1(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ),
    .O(id03902)
  );

  defparam id01753.INIT = 16'h9669;
  LUT4 id01753 (
    .ADR0(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x1 ),
    .ADR2(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR3(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x2 ),
    .O(id03899)
  );

  defparam id01754.INIT = 16'h0D57;
  LUT4 id01754 (
    .ADR0(id03903),
    .ADR1(id03907),
    .ADR2(id03908),
    .ADR3(id03910),
    .O(id03896)
  );

  defparam id01755.INIT = 16'h07F8;
  LUT4 id01755 (
    .ADR0(id03901),
    .ADR1(id03900),
    .ADR2(id03889),
    .ADR3(id03890),
    .O(id03898)
  );

  defparam id01756.INIT = 16'h8700;
  LUT4 id01756 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ),
    .ADR2(id03899),
    .ADR3(id03902),
    .O(id03889)
  );

  defparam id01757.INIT = 4'h9;
  LUT2 id01757 (
    .ADR0(id03887),
    .ADR1(id03888),
    .O(id03890)
  );

  defparam id01758.INIT = 16'h0F77;
  LUT4 id01758 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_0.CELLS[3].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x0 ),
    .ADR3(id03899),
    .O(id03887)
  );

  defparam id01759.INIT = 4'h9;
  LUT2 id01759 (
    .ADR0(id03893),
    .ADR1(id03894),
    .O(id03888)
  );

  defparam id01760.INIT = 16'h9669;
  LUT4 id01760 (
    .ADR0(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x2 ),
    .O(id03893)
  );

  defparam id01761.INIT = 8'hE8;
  LUT3 id01761 (
    .ADR0(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x1 ),
    .ADR1(\DECODE_GEN[2].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_0.CELLS[4].u_compressor42_cell.x2 ),
    .O(id03894)
  );

  defparam id01762.INIT = 4'h8;
  LUT2 id01762 (
    .ADR0(id03908),
    .ADR1(id03910),
    .O(id03900)
  );

  defparam id01763.INIT = 16'h0BF4;
  LUT4 id01763 (
    .ADR0(id03897),
    .ADR1(id03898),
    .ADR2(id03891),
    .ADR3(id03892),
    .O(\net_Buf-pad-result[6] )
  );

  defparam id01764.INIT = 8'h80;
  LUT3 id01764 (
    .ADR0(id03901),
    .ADR1(id03890),
    .ADR2(id03900),
    .O(id03891)
  );

  defparam id01765.INIT = 8'h78;
  LUT3 id01765 (
    .ADR0(id03889),
    .ADR1(id03890),
    .ADR2(id04073),
    .O(id03892)
  );

  defparam id01766.INIT = 16'h4BB4;
  LUT4 id01766 (
    .ADR0(id03887),
    .ADR1(id03888),
    .ADR2(id04074),
    .ADR3(id04071),
    .O(id04073)
  );

  defparam id01767.INIT = 16'h53AC;
  LUT4 id01767 (
    .ADR0(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x0 ),
    .ADR1(id03894),
    .ADR2(id03893),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id04074)
  );

  defparam id01768.INIT = 4'h9;
  LUT2 id01768 (
    .ADR0(id04072),
    .ADR1(id04077),
    .O(id04071)
  );

  defparam id01769.INIT = 16'h9669;
  LUT4 id01769 (
    .ADR0(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04072)
  );

  defparam id01770.INIT = 8'hE8;
  LUT3 id01770 (
    .ADR0(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x1 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x2 ),
    .O(id04077)
  );

  defparam id01771.INIT = 4'h6;
  LUT2 id01771 (
    .ADR0(id04078),
    .ADR1(id04075),
    .O(\net_Buf-pad-result[7] )
  );

  defparam id01772.INIT = 16'hF400;
  LUT4 id01772 (
    .ADR0(id03897),
    .ADR1(id03898),
    .ADR2(id03891),
    .ADR3(id03892),
    .O(id04078)
  );

  defparam id01773.INIT = 4'h6;
  LUT2 id01773 (
    .ADR0(id04076),
    .ADR1(id04065),
    .O(id04075)
  );

  defparam id01774.INIT = 16'h007F;
  LUT4 id01774 (
    .ADR0(id04073),
    .ADR1(id03890),
    .ADR2(id03889),
    .ADR3(id04066),
    .O(id04076)
  );

  defparam id01775.INIT = 16'h1400;
  LUT4 id01775 (
    .ADR0(id03887),
    .ADR1(id04074),
    .ADR2(id04071),
    .ADR3(id03888),
    .O(id04066)
  );

  defparam id01776.INIT = 8'hE1;
  LUT3 id01776 (
    .ADR0(id04063),
    .ADR1(id04064),
    .ADR2(id04069),
    .O(id04065)
  );

  defparam id01777.INIT = 4'h8;
  LUT2 id01777 (
    .ADR0(id04074),
    .ADR1(id04071),
    .O(id04063)
  );

  defparam id01778.INIT = 8'h69;
  LUT3 id01778 (
    .ADR0(id04070),
    .ADR1(id04067),
    .ADR2(GND_NET),
    .O(id04069)
  );

  defparam id01779.INIT = 8'h35;
  LUT3 id01779 (
    .ADR0(id04077),
    .ADR1(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x0 ),
    .ADR2(id04072),
    .O(id04070)
  );

  defparam id01780.INIT = 4'h9;
  LUT2 id01780 (
    .ADR0(id04068),
    .ADR1(id04057),
    .O(id04067)
  );

  defparam id01781.INIT = 16'h9669;
  LUT4 id01781 (
    .ADR0(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04068)
  );

  defparam id01782.INIT = 8'hE8;
  LUT3 id01782 (
    .ADR0(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04057)
  );

  defparam id01783.INIT = 16'hCA00;
  LUT4 id01783 (
    .ADR0(id03894),
    .ADR1(\u_compressor42_l0_0.CELLS[5].u_compressor42_cell.x0 ),
    .ADR2(id03893),
    .ADR3(\DECODE_GEN[3].u_booth_enc.partial_reverse ),
    .O(id04064)
  );

  defparam id01784.INIT = 16'hF807;
  LUT4 id01784 (
    .ADR0(id04078),
    .ADR1(id04075),
    .ADR2(id04058),
    .ADR3(id04055),
    .O(\net_Buf-pad-result[8] )
  );

  defparam id01785.INIT = 16'h4000;
  LUT4 id01785 (
    .ADR0(id04065),
    .ADR1(id03889),
    .ADR2(id03890),
    .ADR3(id04073),
    .O(id04058)
  );

  defparam id01786.INIT = 4'h6;
  LUT2 id01786 (
    .ADR0(id04056),
    .ADR1(id04061),
    .O(id04055)
  );

  defparam id01787.INIT = 4'h6;
  LUT2 id01787 (
    .ADR0(id04062),
    .ADR1(id04059),
    .O(id04056)
  );

  defparam id01788.INIT = 8'h96;
  LUT3 id01788 (
    .ADR0(id04060),
    .ADR1(id04049),
    .ADR2(id04050),
    .O(id04062)
  );

  defparam id01789.INIT = 16'hCA00;
  LUT4 id01789 (
    .ADR0(id04077),
    .ADR1(\u_compressor42_l0_0.CELLS[6].u_compressor42_cell.x0 ),
    .ADR2(id04072),
    .ADR3(GND_NET),
    .O(id04060)
  );

  defparam id01790.INIT = 16'h53AC;
  LUT4 id01790 (
    .ADR0(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x0 ),
    .ADR1(id04057),
    .ADR2(id04068),
    .ADR3(id04047),
    .O(id04049)
  );

  defparam id01791.INIT = 4'h6;
  LUT2 id01791 (
    .ADR0(\u_compressor42_l0_1.CELLS[2].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .O(id04047)
  );

  defparam id01792.INIT = 4'h9;
  LUT2 id01792 (
    .ADR0(id04048),
    .ADR1(id04053),
    .O(id04050)
  );

  defparam id01793.INIT = 16'h9669;
  LUT4 id01793 (
    .ADR0(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04048)
  );

  defparam id01794.INIT = 8'hE8;
  LUT3 id01794 (
    .ADR0(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04053)
  );

  defparam id01795.INIT = 16'hE88E;
  LUT4 id01795 (
    .ADR0(id04064),
    .ADR1(id04067),
    .ADR2(id04070),
    .ADR3(GND_NET),
    .O(id04059)
  );

  defparam id01796.INIT = 16'h0D57;
  LUT4 id01796 (
    .ADR0(id04066),
    .ADR1(id04064),
    .ADR2(id04063),
    .ADR3(id04069),
    .O(id04061)
  );

  defparam id01797.INIT = 8'h1E;
  LUT3 id01797 (
    .ADR0(id04054),
    .ADR1(id04051),
    .ADR2(id04052),
    .O(\net_Buf-pad-result[9] )
  );

  defparam id01798.INIT = 16'h00F8;
  LUT4 id01798 (
    .ADR0(id04075),
    .ADR1(id04078),
    .ADR2(id04058),
    .ADR3(id04055),
    .O(id04054)
  );

  defparam id01799.INIT = 8'h96;
  LUT3 id01799 (
    .ADR0(id04105),
    .ADR1(id04106),
    .ADR2(id04103),
    .O(id04052)
  );

  defparam id01800.INIT = 8'h80;
  LUT3 id01800 (
    .ADR0(id04056),
    .ADR1(id04063),
    .ADR2(id04069),
    .O(id04105)
  );

  defparam id01801.INIT = 4'h8;
  LUT2 id01801 (
    .ADR0(id04062),
    .ADR1(id04059),
    .O(id04106)
  );

  defparam id01802.INIT = 4'h9;
  LUT2 id01802 (
    .ADR0(id04104),
    .ADR1(id04109),
    .O(id04103)
  );

  defparam id01803.INIT = 8'h17;
  LUT3 id01803 (
    .ADR0(id04060),
    .ADR1(id04049),
    .ADR2(id04050),
    .O(id04104)
  );

  defparam id01804.INIT = 16'h9669;
  LUT4 id01804 (
    .ADR0(id04110),
    .ADR1(id04107),
    .ADR2(id04108),
    .ADR3(id04097),
    .O(id04109)
  );

  defparam id01805.INIT = 16'hCA00;
  LUT4 id01805 (
    .ADR0(id04057),
    .ADR1(\u_compressor42_l0_0.CELLS[7].u_compressor42_cell.x0 ),
    .ADR2(id04068),
    .ADR3(id04047),
    .O(id04110)
  );

  defparam id01806.INIT = 4'h9;
  LUT2 id01806 (
    .ADR0(id04098),
    .ADR1(id04095),
    .O(id04107)
  );

  defparam id01807.INIT = 16'h9669;
  LUT4 id01807 (
    .ADR0(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04098)
  );

  defparam id01808.INIT = 8'hE8;
  LUT3 id01808 (
    .ADR0(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04095)
  );

  defparam id01809.INIT = 8'h35;
  LUT3 id01809 (
    .ADR0(id04053),
    .ADR1(\u_compressor42_l0_0.CELLS[8].u_compressor42_cell.x0 ),
    .ADR2(id04048),
    .O(id04108)
  );

  defparam id01810.INIT = 8'h96;
  LUT3 id01810 (
    .ADR0(id04096),
    .ADR1(\u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .O(id04097)
  );

  defparam id01811.INIT = 4'h8;
  LUT2 id01811 (
    .ADR0(\u_compressor42_l0_1.CELLS[2].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[4].u_booth_enc.partial_reverse ),
    .O(id04096)
  );

  defparam id01812.INIT = 8'h40;
  LUT3 id01812 (
    .ADR0(id04065),
    .ADR1(id04056),
    .ADR2(id04066),
    .O(id04051)
  );

  defparam id01813.INIT = 8'h69;
  LUT3 id01813 (
    .ADR0(id04101),
    .ADR1(id04102),
    .ADR2(id04099),
    .O(\net_Buf-pad-result[10] )
  );

  defparam id01814.INIT = 16'h01FF;
  LUT4 id01814 (
    .ADR0(id04051),
    .ADR1(id04105),
    .ADR2(id04054),
    .ADR3(id04103),
    .O(id04101)
  );

  defparam id01815.INIT = 4'h6;
  LUT2 id01815 (
    .ADR0(id04100),
    .ADR1(id04089),
    .O(id04102)
  );

  defparam id01816.INIT = 4'h6;
  LUT2 id01816 (
    .ADR0(id04090),
    .ADR1(id04087),
    .O(id04100)
  );

  defparam id01817.INIT = 8'h96;
  LUT3 id01817 (
    .ADR0(id04088),
    .ADR1(id04093),
    .ADR2(id04094),
    .O(id04090)
  );

  defparam id01818.INIT = 16'h4DD4;
  LUT4 id01818 (
    .ADR0(id04108),
    .ADR1(id04096),
    .ADR2(\u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04088)
  );

  defparam id01819.INIT = 16'h8778;
  LUT4 id01819 (
    .ADR0(\u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(id04091),
    .ADR3(id04092),
    .O(id04093)
  );

  defparam id01820.INIT = 4'h9;
  LUT2 id01820 (
    .ADR0(id04081),
    .ADR1(id04082),
    .O(id04091)
  );

  defparam id01821.INIT = 16'h9669;
  LUT4 id01821 (
    .ADR0(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04081)
  );

  defparam id01822.INIT = 8'hE8;
  LUT3 id01822 (
    .ADR0(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04082)
  );

  defparam id01823.INIT = 8'h96;
  LUT3 id01823 (
    .ADR0(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 ),
    .O(id04092)
  );

  defparam id01824.INIT = 8'h35;
  LUT3 id01824 (
    .ADR0(id04095),
    .ADR1(\u_compressor42_l0_0.CELLS[9].u_compressor42_cell.x0 ),
    .ADR2(id04098),
    .O(id04094)
  );

  defparam id01825.INIT = 16'h1771;
  LUT4 id01825 (
    .ADR0(id04110),
    .ADR1(id04107),
    .ADR2(id04108),
    .ADR3(id04097),
    .O(id04087)
  );

  defparam id01826.INIT = 4'h4;
  LUT2 id01826 (
    .ADR0(id04104),
    .ADR1(id04109),
    .O(id04089)
  );

  defparam id01827.INIT = 4'h8;
  LUT2 id01827 (
    .ADR0(id04106),
    .ADR1(id04103),
    .O(id04099)
  );

  defparam id01828.INIT = 16'hD42B;
  LUT4 id01828 (
    .ADR0(id04101),
    .ADR1(id04102),
    .ADR2(id04099),
    .ADR3(id04079),
    .O(\net_Buf-pad-result[11] )
  );

  defparam id01829.INIT = 8'hE1;
  LUT3 id01829 (
    .ADR0(id04080),
    .ADR1(id04085),
    .ADR2(id04086),
    .O(id04079)
  );

  defparam id01830.INIT = 4'h8;
  LUT2 id01830 (
    .ADR0(id04100),
    .ADR1(id04089),
    .O(id04080)
  );

  defparam id01831.INIT = 4'h1;
  LUT2 id01831 (
    .ADR0(id04090),
    .ADR1(id04087),
    .O(id04085)
  );

  defparam id01832.INIT = 4'h6;
  LUT2 id01832 (
    .ADR0(id04083),
    .ADR1(id04084),
    .O(id04086)
  );

  defparam id01833.INIT = 16'hACCA;
  LUT4 id01833 (
    .ADR0(id04088),
    .ADR1(id04091),
    .ADR2(id04093),
    .ADR3(id04094),
    .O(id04083)
  );

  defparam id01834.INIT = 4'h6;
  LUT2 id01834 (
    .ADR0(id04009),
    .ADR1(id04010),
    .O(id04084)
  );

  defparam id01835.INIT = 16'h1EE1;
  LUT4 id01835 (
    .ADR0(id04007),
    .ADR1(id04008),
    .ADR2(id04013),
    .ADR3(id04014),
    .O(id04009)
  );

  defparam id01836.INIT = 16'h6000;
  LUT4 id01836 (
    .ADR0(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 ),
    .ADR2(id04011),
    .ADR3(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x0 ),
    .O(id04007)
  );

  defparam id01837.INIT = 8'h96;
  LUT3 id01837 (
    .ADR0(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 ),
    .O(id04011)
  );

  defparam id01838.INIT = 16'hC017;
  LUT4 id01838 (
    .ADR0(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 ),
    .ADR3(id04011),
    .O(id04008)
  );

  defparam id01839.INIT = 8'h35;
  LUT3 id01839 (
    .ADR0(id04082),
    .ADR1(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x0 ),
    .ADR2(id04081),
    .O(id04013)
  );

  defparam id01840.INIT = 4'h9;
  LUT2 id01840 (
    .ADR0(id04012),
    .ADR1(id04001),
    .O(id04014)
  );

  defparam id01841.INIT = 16'h9669;
  LUT4 id01841 (
    .ADR0(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x2 ),
    .O(id04012)
  );

  defparam id01842.INIT = 8'hE8;
  LUT3 id01842 (
    .ADR0(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04001)
  );

  defparam id01843.INIT = 16'h2BBB;
  LUT4 id01843 (
    .ADR0(id04094),
    .ADR1(id04092),
    .ADR2(\u_compressor42_l0_1.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04010)
  );

  defparam id01844.INIT = 16'hE11E;
  LUT4 id01844 (
    .ADR0(id04002),
    .ADR1(id03999),
    .ADR2(id04000),
    .ADR3(id04005),
    .O(\net_Buf-pad-result[12] )
  );

  defparam id01845.INIT = 16'h00D4;
  LUT4 id01845 (
    .ADR0(id04101),
    .ADR1(id04102),
    .ADR2(id04099),
    .ADR3(id04079),
    .O(id04002)
  );

  defparam id01846.INIT = 4'h8;
  LUT2 id01846 (
    .ADR0(id04080),
    .ADR1(id04086),
    .O(id03999)
  );

  defparam id01847.INIT = 4'h8;
  LUT2 id01847 (
    .ADR0(id04085),
    .ADR1(id04086),
    .O(id04000)
  );

  defparam id01848.INIT = 4'h6;
  LUT2 id01848 (
    .ADR0(id04006),
    .ADR1(id04003),
    .O(id04005)
  );

  defparam id01849.INIT = 4'h8;
  LUT2 id01849 (
    .ADR0(id04083),
    .ADR1(id04084),
    .O(id04006)
  );

  defparam id01850.INIT = 4'h9;
  LUT2 id01850 (
    .ADR0(id04004),
    .ADR1(id03993),
    .O(id04003)
  );

  defparam id01851.INIT = 8'h3A;
  LUT3 id01851 (
    .ADR0(id04010),
    .ADR1(id04014),
    .ADR2(id04009),
    .O(id04004)
  );

  defparam id01852.INIT = 4'h9;
  LUT2 id01852 (
    .ADR0(id03994),
    .ADR1(id03991),
    .O(id03993)
  );

  defparam id01853.INIT = 16'h9669;
  LUT4 id01853 (
    .ADR0(id03992),
    .ADR1(id03997),
    .ADR2(id03998),
    .ADR3(id03995),
    .O(id03994)
  );

  defparam id01854.INIT = 16'h7117;
  LUT4 id01854 (
    .ADR0(id03996),
    .ADR1(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 ),
    .O(id03992)
  );

  defparam id01855.INIT = 4'h8;
  LUT2 id01855 (
    .ADR0(\DECODE_GEN[5].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_1.CELLS[4].u_compressor42_cell.x1 ),
    .O(id03996)
  );

  defparam id01856.INIT = 8'h87;
  LUT3 id01856 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(id03985),
    .O(id03997)
  );

  defparam id01857.INIT = 16'h9669;
  LUT4 id01857 (
    .ADR0(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x1 ),
    .ADR2(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR3(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x2 ),
    .O(id03985)
  );

  defparam id01858.INIT = 8'h35;
  LUT3 id01858 (
    .ADR0(id04001),
    .ADR1(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x0 ),
    .ADR2(id04012),
    .O(id03998)
  );

  defparam id01859.INIT = 4'h9;
  LUT2 id01859 (
    .ADR0(id03986),
    .ADR1(id03983),
    .O(id03995)
  );

  defparam id01860.INIT = 16'h9669;
  LUT4 id01860 (
    .ADR0(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x2 ),
    .O(id03986)
  );

  defparam id01861.INIT = 8'hE8;
  LUT3 id01861 (
    .ADR0(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[11].u_compressor42_cell.x2 ),
    .O(id03983)
  );

  defparam id01862.INIT = 8'h0D;
  LUT3 id01862 (
    .ADR0(id04013),
    .ADR1(id04007),
    .ADR2(id04008),
    .O(id03991)
  );

  defparam id01863.INIT = 4'h9;
  LUT2 id01863 (
    .ADR0(id03984),
    .ADR1(id03989),
    .O(\net_Buf-pad-result[13] )
  );

  defparam id01864.INIT = 16'h1117;
  LUT4 id01864 (
    .ADR0(id04000),
    .ADR1(id04005),
    .ADR2(id04002),
    .ADR3(id03999),
    .O(id03984)
  );

  defparam id01865.INIT = 8'h1E;
  LUT3 id01865 (
    .ADR0(id03990),
    .ADR1(id03987),
    .ADR2(id03988),
    .O(id03989)
  );

  defparam id01866.INIT = 4'h8;
  LUT2 id01866 (
    .ADR0(id04006),
    .ADR1(id04003),
    .O(id03990)
  );

  defparam id01867.INIT = 4'h4;
  LUT2 id01867 (
    .ADR0(id04004),
    .ADR1(id03993),
    .O(id03987)
  );

  defparam id01868.INIT = 4'h9;
  LUT2 id01868 (
    .ADR0(id04041),
    .ADR1(id04042),
    .O(id03988)
  );

  defparam id01869.INIT = 8'h35;
  LUT3 id01869 (
    .ADR0(id03991),
    .ADR1(id03995),
    .ADR2(id03994),
    .O(id04041)
  );

  defparam id01870.INIT = 4'h9;
  LUT2 id01870 (
    .ADR0(id04039),
    .ADR1(id04040),
    .O(id04042)
  );

  defparam id01871.INIT = 16'h6996;
  LUT4 id01871 (
    .ADR0(id04045),
    .ADR1(id04046),
    .ADR2(id04043),
    .ADR3(id04044),
    .O(id04039)
  );

  defparam id01872.INIT = 16'h0F77;
  LUT4 id01872 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_1.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x0 ),
    .ADR3(id03985),
    .O(id04045)
  );

  defparam id01873.INIT = 4'h9;
  LUT2 id01873 (
    .ADR0(id04033),
    .ADR1(id04034),
    .O(id04046)
  );

  defparam id01874.INIT = 16'h9669;
  LUT4 id01874 (
    .ADR0(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x1 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04033)
  );

  defparam id01875.INIT = 8'hE8;
  LUT3 id01875 (
    .ADR0(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x1 ),
    .ADR1(\DECODE_GEN[6].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_1.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04034)
  );

  defparam id01876.INIT = 8'h35;
  LUT3 id01876 (
    .ADR0(id03983),
    .ADR1(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x0 ),
    .ADR2(id03986),
    .O(id04043)
  );

  defparam id01877.INIT = 4'h9;
  LUT2 id01877 (
    .ADR0(id04031),
    .ADR1(id04032),
    .O(id04044)
  );

  defparam id01878.INIT = 16'h9669;
  LUT4 id01878 (
    .ADR0(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04031)
  );

  defparam id01879.INIT = 8'hE8;
  LUT3 id01879 (
    .ADR0(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[12].u_compressor42_cell.x2 ),
    .O(id04032)
  );

  defparam id01880.INIT = 8'hB2;
  LUT3 id01880 (
    .ADR0(id03992),
    .ADR1(id03997),
    .ADR2(id03998),
    .O(id04040)
  );

  defparam id01881.INIT = 16'h0BF4;
  LUT4 id01881 (
    .ADR0(id03984),
    .ADR1(id03989),
    .ADR2(id04037),
    .ADR3(id04038),
    .O(\net_Buf-pad-result[14] )
  );

  defparam id01882.INIT = 4'h8;
  LUT2 id01882 (
    .ADR0(id03990),
    .ADR1(id03988),
    .O(id04037)
  );

  defparam id01883.INIT = 8'h1E;
  LUT3 id01883 (
    .ADR0(id04035),
    .ADR1(id04036),
    .ADR2(id04025),
    .O(id04038)
  );

  defparam id01884.INIT = 4'h8;
  LUT2 id01884 (
    .ADR0(id03987),
    .ADR1(id03988),
    .O(id04035)
  );

  defparam id01885.INIT = 4'h6;
  LUT2 id01885 (
    .ADR0(id04026),
    .ADR1(id04023),
    .O(id04025)
  );

  defparam id01886.INIT = 4'h9;
  LUT2 id01886 (
    .ADR0(id04024),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .O(id04026)
  );

  defparam id01887.INIT = 8'hC5;
  LUT3 id01887 (
    .ADR0(id04044),
    .ADR1(id04040),
    .ADR2(id04039),
    .O(id04024)
  );

  defparam id01888.INIT = 4'h6;
  LUT2 id01888 (
    .ADR0(id04029),
    .ADR1(id04030),
    .O(id04023)
  );

  defparam id01889.INIT = 16'h9669;
  LUT4 id01889 (
    .ADR0(id04027),
    .ADR1(id04028),
    .ADR2(id04017),
    .ADR3(id04018),
    .O(id04029)
  );

  defparam id01890.INIT = 8'h35;
  LUT3 id01890 (
    .ADR0(id04034),
    .ADR1(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x0 ),
    .ADR2(id04033),
    .O(id04027)
  );

  defparam id01891.INIT = 4'h9;
  LUT2 id01891 (
    .ADR0(id04015),
    .ADR1(id04016),
    .O(id04028)
  );

  defparam id01892.INIT = 16'h9669;
  LUT4 id01892 (
    .ADR0(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04015)
  );

  defparam id01893.INIT = 8'hE8;
  LUT3 id01893 (
    .ADR0(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x1 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_1.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04016)
  );

  defparam id01894.INIT = 8'h35;
  LUT3 id01894 (
    .ADR0(id04032),
    .ADR1(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x0 ),
    .ADR2(id04031),
    .O(id04017)
  );

  defparam id01895.INIT = 4'h9;
  LUT2 id01895 (
    .ADR0(id04021),
    .ADR1(id04022),
    .O(id04018)
  );

  defparam id01896.INIT = 16'h9669;
  LUT4 id01896 (
    .ADR0(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04021)
  );

  defparam id01897.INIT = 8'hE8;
  LUT3 id01897 (
    .ADR0(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04022)
  );

  defparam id01898.INIT = 8'hB2;
  LUT3 id01898 (
    .ADR0(id04045),
    .ADR1(id04046),
    .ADR2(id04043),
    .O(id04030)
  );

  defparam id01899.INIT = 4'h4;
  LUT2 id01899 (
    .ADR0(id04041),
    .ADR1(id04042),
    .O(id04036)
  );

  defparam id01900.INIT = 8'h1E;
  LUT3 id01900 (
    .ADR0(id04019),
    .ADR1(id04020),
    .ADR2(id04201),
    .O(\net_Buf-pad-result[15] )
  );

  defparam id01901.INIT = 16'hF400;
  LUT4 id01901 (
    .ADR0(id03984),
    .ADR1(id03989),
    .ADR2(id04037),
    .ADR3(id04038),
    .O(id04019)
  );

  defparam id01902.INIT = 8'h1E;
  LUT3 id01902 (
    .ADR0(id04202),
    .ADR1(id04199),
    .ADR2(id04200),
    .O(id04201)
  );

  defparam id01903.INIT = 4'h8;
  LUT2 id01903 (
    .ADR0(id04025),
    .ADR1(id04036),
    .O(id04202)
  );

  defparam id01904.INIT = 4'h8;
  LUT2 id01904 (
    .ADR0(id04026),
    .ADR1(id04023),
    .O(id04199)
  );

  defparam id01905.INIT = 8'h96;
  LUT3 id01905 (
    .ADR0(id04205),
    .ADR1(id04206),
    .ADR2(id04203),
    .O(id04200)
  );

  defparam id01906.INIT = 4'h4;
  LUT2 id01906 (
    .ADR0(id04024),
    .ADR1(\DECODE_GEN[7].u_booth_enc.partial_reverse ),
    .O(id04205)
  );

  defparam id01907.INIT = 4'h9;
  LUT2 id01907 (
    .ADR0(id04204),
    .ADR1(GND_NET),
    .O(id04206)
  );

  defparam id01908.INIT = 8'h3A;
  LUT3 id01908 (
    .ADR0(id04030),
    .ADR1(id04018),
    .ADR2(id04029),
    .O(id04204)
  );

  defparam id01909.INIT = 4'h6;
  LUT2 id01909 (
    .ADR0(id04193),
    .ADR1(id04194),
    .O(id04203)
  );

  defparam id01910.INIT = 16'h9669;
  LUT4 id01910 (
    .ADR0(id04191),
    .ADR1(id04192),
    .ADR2(id04197),
    .ADR3(id04198),
    .O(id04193)
  );

  defparam id01911.INIT = 8'h35;
  LUT3 id01911 (
    .ADR0(id04016),
    .ADR1(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x0 ),
    .ADR2(id04015),
    .O(id04191)
  );

  defparam id01912.INIT = 4'h9;
  LUT2 id01912 (
    .ADR0(id04195),
    .ADR1(id04196),
    .O(id04192)
  );

  defparam id01913.INIT = 16'h9669;
  LUT4 id01913 (
    .ADR0(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04195)
  );

  defparam id01914.INIT = 8'hE8;
  LUT3 id01914 (
    .ADR0(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04196)
  );

  defparam id01915.INIT = 8'h35;
  LUT3 id01915 (
    .ADR0(id04022),
    .ADR1(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x0 ),
    .ADR2(id04021),
    .O(id04197)
  );

  defparam id01916.INIT = 16'h6996;
  LUT4 id01916 (
    .ADR0(id04185),
    .ADR1(id04186),
    .ADR2(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x3 ),
    .O(id04198)
  );

  defparam id01917.INIT = 4'h6;
  LUT2 id01917 (
    .ADR0(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04185)
  );

  defparam id01918.INIT = 8'hE8;
  LUT3 id01918 (
    .ADR0(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04186)
  );

  defparam id01919.INIT = 8'hB2;
  LUT3 id01919 (
    .ADR0(id04027),
    .ADR1(id04028),
    .ADR2(id04017),
    .O(id04194)
  );

  defparam id01920.INIT = 4'h8;
  LUT2 id01920 (
    .ADR0(id04035),
    .ADR1(id04025),
    .O(id04020)
  );

  defparam id01921.INIT = 4'h9;
  LUT2 id01921 (
    .ADR0(id04183),
    .ADR1(id04184),
    .O(\net_Buf-pad-result[16] )
  );

  defparam id01922.INIT = 16'h03FD;
  LUT4 id01922 (
    .ADR0(id04202),
    .ADR1(id04019),
    .ADR2(id04020),
    .ADR3(id04201),
    .O(id04183)
  );

  defparam id01923.INIT = 4'h6;
  LUT2 id01923 (
    .ADR0(id04189),
    .ADR1(id04190),
    .O(id04184)
  );

  defparam id01924.INIT = 4'h8;
  LUT2 id01924 (
    .ADR0(id04199),
    .ADR1(id04200),
    .O(id04189)
  );

  defparam id01925.INIT = 4'h9;
  LUT2 id01925 (
    .ADR0(id04187),
    .ADR1(id04188),
    .O(id04190)
  );

  defparam id01926.INIT = 8'h17;
  LUT3 id01926 (
    .ADR0(id04205),
    .ADR1(id04206),
    .ADR2(id04203),
    .O(id04187)
  );

  defparam id01927.INIT = 8'h96;
  LUT3 id01927 (
    .ADR0(id04177),
    .ADR1(id04178),
    .ADR2(id04175),
    .O(id04188)
  );

  defparam id01928.INIT = 4'h4;
  LUT2 id01928 (
    .ADR0(id04204),
    .ADR1(GND_NET),
    .O(id04177)
  );

  defparam id01929.INIT = 8'h69;
  LUT3 id01929 (
    .ADR0(id04176),
    .ADR1(\u_compressor42_l0_2.CELLS[2].u_compressor42_cell.x0 ),
    .ADR2(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .O(id04178)
  );

  defparam id01930.INIT = 8'h3A;
  LUT3 id01930 (
    .ADR0(id04194),
    .ADR1(id04198),
    .ADR2(id04193),
    .O(id04176)
  );

  defparam id01931.INIT = 4'h9;
  LUT2 id01931 (
    .ADR0(id04181),
    .ADR1(id04182),
    .O(id04175)
  );

  defparam id01932.INIT = 16'h6996;
  LUT4 id01932 (
    .ADR0(id04179),
    .ADR1(id04180),
    .ADR2(id04233),
    .ADR3(id04234),
    .O(id04181)
  );

  defparam id01933.INIT = 8'h35;
  LUT3 id01933 (
    .ADR0(id04196),
    .ADR1(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x0 ),
    .ADR2(id04195),
    .O(id04179)
  );

  defparam id01934.INIT = 4'h9;
  LUT2 id01934 (
    .ADR0(id04231),
    .ADR1(id04232),
    .O(id04180)
  );

  defparam id01935.INIT = 16'h9669;
  LUT4 id01935 (
    .ADR0(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04231)
  );

  defparam id01936.INIT = 8'hE8;
  LUT3 id01936 (
    .ADR0(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04232)
  );

  defparam id01937.INIT = 16'h7117;
  LUT4 id01937 (
    .ADR0(id04186),
    .ADR1(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x0 ),
    .ADR2(id04185),
    .ADR3(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x3 ),
    .O(id04233)
  );

  defparam id01938.INIT = 4'h9;
  LUT2 id01938 (
    .ADR0(id04237),
    .ADR1(id04238),
    .O(id04234)
  );

  defparam id01939.INIT = 16'h9669;
  LUT4 id01939 (
    .ADR0(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04237)
  );

  defparam id01940.INIT = 8'hE8;
  LUT3 id01940 (
    .ADR0(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04238)
  );

  defparam id01941.INIT = 8'hB2;
  LUT3 id01941 (
    .ADR0(id04191),
    .ADR1(id04192),
    .ADR2(id04197),
    .O(id04182)
  );

  defparam id01942.INIT = 16'h2BD4;
  LUT4 id01942 (
    .ADR0(id04183),
    .ADR1(id04189),
    .ADR2(id04190),
    .ADR3(id04235),
    .O(\net_Buf-pad-result[17] )
  );

  defparam id01943.INIT = 4'h6;
  LUT2 id01943 (
    .ADR0(id04236),
    .ADR1(id04225),
    .O(id04235)
  );

  defparam id01944.INIT = 4'h4;
  LUT2 id01944 (
    .ADR0(id04187),
    .ADR1(id04188),
    .O(id04236)
  );

  defparam id01945.INIT = 4'h9;
  LUT2 id01945 (
    .ADR0(id04226),
    .ADR1(id04223),
    .O(id04225)
  );

  defparam id01946.INIT = 8'h17;
  LUT3 id01946 (
    .ADR0(id04177),
    .ADR1(id04178),
    .ADR2(id04175),
    .O(id04226)
  );

  defparam id01947.INIT = 8'h96;
  LUT3 id01947 (
    .ADR0(id04224),
    .ADR1(id04229),
    .ADR2(id04230),
    .O(id04223)
  );

  defparam id01948.INIT = 8'h14;
  LUT3 id01948 (
    .ADR0(id04176),
    .ADR1(\u_compressor42_l0_2.CELLS[2].u_compressor42_cell.x0 ),
    .ADR2(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .O(id04224)
  );

  defparam id01949.INIT = 16'h9669;
  LUT4 id01949 (
    .ADR0(id04227),
    .ADR1(id04228),
    .ADR2(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04229)
  );

  defparam id01950.INIT = 8'hC5;
  LUT3 id01950 (
    .ADR0(id04234),
    .ADR1(id04182),
    .ADR2(id04181),
    .O(id04227)
  );

  defparam id01951.INIT = 4'h8;
  LUT2 id01951 (
    .ADR0(\u_compressor42_l0_2.CELLS[2].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[8].u_booth_enc.partial_reverse ),
    .O(id04228)
  );

  defparam id01952.INIT = 4'h9;
  LUT2 id01952 (
    .ADR0(id04217),
    .ADR1(id04218),
    .O(id04230)
  );

  defparam id01953.INIT = 16'h6996;
  LUT4 id01953 (
    .ADR0(id04215),
    .ADR1(id04216),
    .ADR2(id04221),
    .ADR3(id04222),
    .O(id04217)
  );

  defparam id01954.INIT = 8'h35;
  LUT3 id01954 (
    .ADR0(id04232),
    .ADR1(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x0 ),
    .ADR2(id04231),
    .O(id04215)
  );

  defparam id01955.INIT = 4'h9;
  LUT2 id01955 (
    .ADR0(id04219),
    .ADR1(id04220),
    .O(id04216)
  );

  defparam id01956.INIT = 16'h9669;
  LUT4 id01956 (
    .ADR0(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x2 ),
    .O(id04219)
  );

  defparam id01957.INIT = 8'hE8;
  LUT3 id01957 (
    .ADR0(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04220)
  );

  defparam id01958.INIT = 8'h35;
  LUT3 id01958 (
    .ADR0(id04238),
    .ADR1(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x0 ),
    .ADR2(id04237),
    .O(id04221)
  );

  defparam id01959.INIT = 16'h6996;
  LUT4 id01959 (
    .ADR0(id04209),
    .ADR1(id04210),
    .ADR2(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x3 ),
    .O(id04222)
  );

  defparam id01960.INIT = 4'h6;
  LUT2 id01960 (
    .ADR0(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04209)
  );

  defparam id01961.INIT = 8'hE8;
  LUT3 id01961 (
    .ADR0(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04210)
  );

  defparam id01962.INIT = 8'hB2;
  LUT3 id01962 (
    .ADR0(id04179),
    .ADR1(id04180),
    .ADR2(id04233),
    .O(id04218)
  );

  defparam id01963.INIT = 4'h9;
  LUT2 id01963 (
    .ADR0(id04207),
    .ADR1(id04208),
    .O(\net_Buf-pad-result[18] )
  );

  defparam id01964.INIT = 16'hBF00;
  LUT4 id01964 (
    .ADR0(id04183),
    .ADR1(id04235),
    .ADR2(id04184),
    .ADR3(id04213),
    .O(id04207)
  );

  defparam id01965.INIT = 16'h1777;
  LUT4 id01965 (
    .ADR0(id04236),
    .ADR1(id04225),
    .ADR2(id04190),
    .ADR3(id04189),
    .O(id04213)
  );

  defparam id01966.INIT = 4'h6;
  LUT2 id01966 (
    .ADR0(id04214),
    .ADR1(id04211),
    .O(id04208)
  );

  defparam id01967.INIT = 4'h4;
  LUT2 id01967 (
    .ADR0(id04226),
    .ADR1(id04223),
    .O(id04214)
  );

  defparam id01968.INIT = 4'h9;
  LUT2 id01968 (
    .ADR0(id04212),
    .ADR1(id04137),
    .O(id04211)
  );

  defparam id01969.INIT = 8'h17;
  LUT3 id01969 (
    .ADR0(id04224),
    .ADR1(id04229),
    .ADR2(id04230),
    .O(id04212)
  );

  defparam id01970.INIT = 4'h9;
  LUT2 id01970 (
    .ADR0(id04138),
    .ADR1(id04135),
    .O(id04137)
  );

  defparam id01971.INIT = 16'h4114;
  LUT4 id01971 (
    .ADR0(id04227),
    .ADR1(id04228),
    .ADR2(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04138)
  );

  defparam id01972.INIT = 16'h1EE1;
  LUT4 id01972 (
    .ADR0(id04136),
    .ADR1(id04141),
    .ADR2(id04142),
    .ADR3(id04139),
    .O(id04135)
  );

  defparam id01973.INIT = 8'hC5;
  LUT3 id01973 (
    .ADR0(id04222),
    .ADR1(id04218),
    .ADR2(id04217),
    .O(id04142)
  );

  defparam id01974.INIT = 4'h6;
  LUT2 id01974 (
    .ADR0(id04140),
    .ADR1(id04129),
    .O(id04139)
  );

  defparam id01975.INIT = 16'h9669;
  LUT4 id01975 (
    .ADR0(id04130),
    .ADR1(id04127),
    .ADR2(id04128),
    .ADR3(id04133),
    .O(id04140)
  );

  defparam id01976.INIT = 8'h35;
  LUT3 id01976 (
    .ADR0(id04220),
    .ADR1(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x0 ),
    .ADR2(id04219),
    .O(id04130)
  );

  defparam id01977.INIT = 4'h9;
  LUT2 id01977 (
    .ADR0(id04134),
    .ADR1(id04131),
    .O(id04127)
  );

  defparam id01978.INIT = 16'h9669;
  LUT4 id01978 (
    .ADR0(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x2 ),
    .O(id04134)
  );

  defparam id01979.INIT = 8'hE8;
  LUT3 id01979 (
    .ADR0(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[11].u_compressor42_cell.x2 ),
    .O(id04131)
  );

  defparam id01980.INIT = 16'h7117;
  LUT4 id01980 (
    .ADR0(id04210),
    .ADR1(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x0 ),
    .ADR2(id04209),
    .ADR3(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x3 ),
    .O(id04128)
  );

  defparam id01981.INIT = 16'h6996;
  LUT4 id01981 (
    .ADR0(id04132),
    .ADR1(id04121),
    .ADR2(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x3 ),
    .O(id04133)
  );

  defparam id01982.INIT = 4'h6;
  LUT2 id01982 (
    .ADR0(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x2 ),
    .O(id04132)
  );

  defparam id01983.INIT = 8'hE8;
  LUT3 id01983 (
    .ADR0(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04121)
  );

  defparam id01984.INIT = 8'hB2;
  LUT3 id01984 (
    .ADR0(id04215),
    .ADR1(id04216),
    .ADR2(id04221),
    .O(id04129)
  );

  defparam id01985.INIT = 16'h6000;
  LUT4 id01985 (
    .ADR0(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(id04228),
    .ADR3(id04122),
    .O(id04136)
  );

  defparam id01986.INIT = 8'h96;
  LUT3 id01986 (
    .ADR0(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x1 ),
    .O(id04122)
  );

  defparam id01987.INIT = 16'hC017;
  LUT4 id01987 (
    .ADR0(id04228),
    .ADR1(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .ADR3(id04122),
    .O(id04141)
  );

  defparam id01988.INIT = 16'h0BF4;
  LUT4 id01988 (
    .ADR0(id04207),
    .ADR1(id04208),
    .ADR2(id04119),
    .ADR3(id04120),
    .O(\net_Buf-pad-result[19] )
  );

  defparam id01989.INIT = 4'h8;
  LUT2 id01989 (
    .ADR0(id04214),
    .ADR1(id04211),
    .O(id04119)
  );

  defparam id01990.INIT = 4'h6;
  LUT2 id01990 (
    .ADR0(id04125),
    .ADR1(id04126),
    .O(id04120)
  );

  defparam id01991.INIT = 4'h4;
  LUT2 id01991 (
    .ADR0(id04212),
    .ADR1(id04137),
    .O(id04125)
  );

  defparam id01992.INIT = 4'h9;
  LUT2 id01992 (
    .ADR0(id04123),
    .ADR1(id04124),
    .O(id04126)
  );

  defparam id01993.INIT = 8'h53;
  LUT3 id01993 (
    .ADR0(id04139),
    .ADR1(id04138),
    .ADR2(id04135),
    .O(id04123)
  );

  defparam id01994.INIT = 8'h96;
  LUT3 id01994 (
    .ADR0(id04113),
    .ADR1(id04114),
    .ADR2(id04111),
    .O(id04124)
  );

  defparam id01995.INIT = 16'h9669;
  LUT4 id01995 (
    .ADR0(id04112),
    .ADR1(id04117),
    .ADR2(id04118),
    .ADR3(id04115),
    .O(id04113)
  );

  defparam id01996.INIT = 8'h3A;
  LUT3 id01996 (
    .ADR0(id04129),
    .ADR1(id04133),
    .ADR2(id04140),
    .O(id04112)
  );

  defparam id01997.INIT = 8'h80;
  LUT3 id01997 (
    .ADR0(id04122),
    .ADR1(\u_compressor42_l0_2.CELLS[3].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .O(id04117)
  );

  defparam id01998.INIT = 4'h1;
  LUT2 id01998 (
    .ADR0(id04116),
    .ADR1(id04169),
    .O(id04118)
  );

  defparam id01999.INIT = 4'h8;
  LUT2 id01999 (
    .ADR0(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x1 ),
    .O(id04116)
  );

  defparam id02000.INIT = 8'h60;
  LUT3 id02000 (
    .ADR0(\DECODE_GEN[9].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_2.CELLS[4].u_compressor42_cell.x0 ),
    .O(id04169)
  );

  defparam id02001.INIT = 8'h96;
  LUT3 id02001 (
    .ADR0(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ),
    .O(id04115)
  );

  defparam id02002.INIT = 8'h0E;
  LUT3 id02002 (
    .ADR0(id04141),
    .ADR1(id04142),
    .ADR2(id04136),
    .O(id04114)
  );

  defparam id02003.INIT = 4'h9;
  LUT2 id02003 (
    .ADR0(id04170),
    .ADR1(id04167),
    .O(id04111)
  );

  defparam id02004.INIT = 16'h6996;
  LUT4 id02004 (
    .ADR0(id04168),
    .ADR1(id04173),
    .ADR2(id04174),
    .ADR3(id04171),
    .O(id04170)
  );

  defparam id02005.INIT = 8'h35;
  LUT3 id02005 (
    .ADR0(id04131),
    .ADR1(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x0 ),
    .ADR2(id04134),
    .O(id04168)
  );

  defparam id02006.INIT = 4'h9;
  LUT2 id02006 (
    .ADR0(id04172),
    .ADR1(id04161),
    .O(id04173)
  );

  defparam id02007.INIT = 16'h9669;
  LUT4 id02007 (
    .ADR0(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04172)
  );

  defparam id02008.INIT = 8'hE8;
  LUT3 id02008 (
    .ADR0(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[12].u_compressor42_cell.x2 ),
    .O(id04161)
  );

  defparam id02009.INIT = 16'h7117;
  LUT4 id02009 (
    .ADR0(id04121),
    .ADR1(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x0 ),
    .ADR2(id04132),
    .ADR3(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x3 ),
    .O(id04174)
  );

  defparam id02010.INIT = 16'h6996;
  LUT4 id02010 (
    .ADR0(id04162),
    .ADR1(id04159),
    .ADR2(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x3 ),
    .O(id04171)
  );

  defparam id02011.INIT = 4'h6;
  LUT2 id02011 (
    .ADR0(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x2 ),
    .O(id04162)
  );

  defparam id02012.INIT = 8'hE8;
  LUT3 id02012 (
    .ADR0(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[18].u_compressor42_cell.x2 ),
    .O(id04159)
  );

  defparam id02013.INIT = 8'hB2;
  LUT3 id02013 (
    .ADR0(id04130),
    .ADR1(id04127),
    .ADR2(id04128),
    .O(id04167)
  );

  defparam id02014.INIT = 4'h9;
  LUT2 id02014 (
    .ADR0(id04160),
    .ADR1(id04165),
    .O(\net_Buf-pad-result[20] )
  );

  defparam id02015.INIT = 16'hBF00;
  LUT4 id02015 (
    .ADR0(id04207),
    .ADR1(id04208),
    .ADR2(id04120),
    .ADR3(id04166),
    .O(id04160)
  );

  defparam id02016.INIT = 8'h1F;
  LUT3 id02016 (
    .ADR0(id04125),
    .ADR1(id04119),
    .ADR2(id04126),
    .O(id04166)
  );

  defparam id02017.INIT = 4'h6;
  LUT2 id02017 (
    .ADR0(id04163),
    .ADR1(id04164),
    .O(id04165)
  );

  defparam id02018.INIT = 4'h4;
  LUT2 id02018 (
    .ADR0(id04123),
    .ADR1(id04124),
    .O(id04163)
  );

  defparam id02019.INIT = 4'h9;
  LUT2 id02019 (
    .ADR0(id04153),
    .ADR1(id04154),
    .O(id04164)
  );

  defparam id02020.INIT = 8'hB2;
  LUT3 id02020 (
    .ADR0(id04113),
    .ADR1(id04111),
    .ADR2(id04114),
    .O(id04153)
  );

  defparam id02021.INIT = 8'h96;
  LUT3 id02021 (
    .ADR0(id04151),
    .ADR1(id04152),
    .ADR2(id04157),
    .O(id04154)
  );

  defparam id02022.INIT = 16'h8778;
  LUT4 id02022 (
    .ADR0(id04169),
    .ADR1(id04115),
    .ADR2(id04158),
    .ADR3(id04155),
    .O(id04151)
  );

  defparam id02023.INIT = 8'hC5;
  LUT3 id02023 (
    .ADR0(id04171),
    .ADR1(id04167),
    .ADR2(id04170),
    .O(id04158)
  );

  defparam id02024.INIT = 16'h7887;
  LUT4 id02024 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(id04156),
    .ADR3(id04145),
    .O(id04155)
  );

  defparam id02025.INIT = 16'h8EE8;
  LUT4 id02025 (
    .ADR0(id04116),
    .ADR1(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ),
    .O(id04156)
  );

  defparam id02026.INIT = 16'h9669;
  LUT4 id02026 (
    .ADR0(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x1 ),
    .ADR2(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR3(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04145)
  );

  defparam id02027.INIT = 16'h2BB2;
  LUT4 id02027 (
    .ADR0(id04112),
    .ADR1(id04117),
    .ADR2(id04118),
    .ADR3(id04115),
    .O(id04152)
  );

  defparam id02028.INIT = 4'h9;
  LUT2 id02028 (
    .ADR0(id04146),
    .ADR1(id04143),
    .O(id04157)
  );

  defparam id02029.INIT = 16'h6996;
  LUT4 id02029 (
    .ADR0(id04144),
    .ADR1(id04149),
    .ADR2(id04150),
    .ADR3(id04147),
    .O(id04146)
  );

  defparam id02030.INIT = 8'h35;
  LUT3 id02030 (
    .ADR0(id04161),
    .ADR1(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x0 ),
    .ADR2(id04172),
    .O(id04144)
  );

  defparam id02031.INIT = 4'h9;
  LUT2 id02031 (
    .ADR0(id04148),
    .ADR1(id04579),
    .O(id04149)
  );

  defparam id02032.INIT = 16'h9669;
  LUT4 id02032 (
    .ADR0(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04148)
  );

  defparam id02033.INIT = 8'hE8;
  LUT3 id02033 (
    .ADR0(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04579)
  );

  defparam id02034.INIT = 16'h7117;
  LUT4 id02034 (
    .ADR0(id04159),
    .ADR1(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x0 ),
    .ADR2(id04162),
    .ADR3(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x3 ),
    .O(id04150)
  );

  defparam id02035.INIT = 16'h6996;
  LUT4 id02035 (
    .ADR0(id04580),
    .ADR1(id04577),
    .ADR2(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x3 ),
    .O(id04147)
  );

  defparam id02036.INIT = 4'h6;
  LUT2 id02036 (
    .ADR0(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x2 ),
    .O(id04580)
  );

  defparam id02037.INIT = 8'hE8;
  LUT3 id02037 (
    .ADR0(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[19].u_compressor42_cell.x2 ),
    .O(id04577)
  );

  defparam id02038.INIT = 8'hB2;
  LUT3 id02038 (
    .ADR0(id04168),
    .ADR1(id04173),
    .ADR2(id04174),
    .O(id04143)
  );

  defparam id02039.INIT = 16'h0BF4;
  LUT4 id02039 (
    .ADR0(id04160),
    .ADR1(id04165),
    .ADR2(id04578),
    .ADR3(id04583),
    .O(\net_Buf-pad-result[21] )
  );

  defparam id02040.INIT = 4'h8;
  LUT2 id02040 (
    .ADR0(id04163),
    .ADR1(id04164),
    .O(id04578)
  );

  defparam id02041.INIT = 4'h6;
  LUT2 id02041 (
    .ADR0(id04584),
    .ADR1(id04581),
    .O(id04583)
  );

  defparam id02042.INIT = 4'h4;
  LUT2 id02042 (
    .ADR0(id04153),
    .ADR1(id04154),
    .O(id04584)
  );

  defparam id02043.INIT = 4'h9;
  LUT2 id02043 (
    .ADR0(id04582),
    .ADR1(id04571),
    .O(id04581)
  );

  defparam id02044.INIT = 8'hB2;
  LUT3 id02044 (
    .ADR0(id04151),
    .ADR1(id04157),
    .ADR2(id04152),
    .O(id04582)
  );

  defparam id02045.INIT = 8'h96;
  LUT3 id02045 (
    .ADR0(id04572),
    .ADR1(id04569),
    .ADR2(id04570),
    .O(id04571)
  );

  defparam id02046.INIT = 8'h96;
  LUT3 id02046 (
    .ADR0(id04575),
    .ADR1(id04576),
    .ADR2(id04573),
    .O(id04572)
  );

  defparam id02047.INIT = 8'hC5;
  LUT3 id02047 (
    .ADR0(id04147),
    .ADR1(id04143),
    .ADR2(id04146),
    .O(id04575)
  );

  defparam id02048.INIT = 16'h8700;
  LUT4 id02048 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(id04145),
    .ADR3(id04156),
    .O(id04576)
  );

  defparam id02049.INIT = 4'h9;
  LUT2 id02049 (
    .ADR0(id04574),
    .ADR1(id04563),
    .O(id04573)
  );

  defparam id02050.INIT = 16'h0F77;
  LUT4 id02050 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_2.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x0 ),
    .ADR3(id04145),
    .O(id04574)
  );

  defparam id02051.INIT = 4'h9;
  LUT2 id02051 (
    .ADR0(id04564),
    .ADR1(id04561),
    .O(id04563)
  );

  defparam id02052.INIT = 16'h9669;
  LUT4 id02052 (
    .ADR0(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x1 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04564)
  );

  defparam id02053.INIT = 8'hE8;
  LUT3 id02053 (
    .ADR0(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x1 ),
    .ADR1(\DECODE_GEN[10].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_2.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04561)
  );

  defparam id02054.INIT = 16'h2BBB;
  LUT4 id02054 (
    .ADR0(id04158),
    .ADR1(id04155),
    .ADR2(id04169),
    .ADR3(id04115),
    .O(id04569)
  );

  defparam id02055.INIT = 4'h9;
  LUT2 id02055 (
    .ADR0(id04562),
    .ADR1(id04567),
    .O(id04570)
  );

  defparam id02056.INIT = 16'h6996;
  LUT4 id02056 (
    .ADR0(id04568),
    .ADR1(id04565),
    .ADR2(id04566),
    .ADR3(id04555),
    .O(id04562)
  );

  defparam id02057.INIT = 8'h35;
  LUT3 id02057 (
    .ADR0(id04579),
    .ADR1(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x0 ),
    .ADR2(id04148),
    .O(id04568)
  );

  defparam id02058.INIT = 4'h9;
  LUT2 id02058 (
    .ADR0(id04556),
    .ADR1(id04553),
    .O(id04565)
  );

  defparam id02059.INIT = 16'h9669;
  LUT4 id02059 (
    .ADR0(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04556)
  );

  defparam id02060.INIT = 8'hE8;
  LUT3 id02060 (
    .ADR0(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04553)
  );

  defparam id02061.INIT = 16'h7117;
  LUT4 id02061 (
    .ADR0(id04577),
    .ADR1(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x0 ),
    .ADR2(id04580),
    .ADR3(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x3 ),
    .O(id04566)
  );

  defparam id02062.INIT = 16'h6996;
  LUT4 id02062 (
    .ADR0(id04554),
    .ADR1(id04559),
    .ADR2(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x3 ),
    .O(id04555)
  );

  defparam id02063.INIT = 4'h6;
  LUT2 id02063 (
    .ADR0(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x2 ),
    .O(id04554)
  );

  defparam id02064.INIT = 8'hE8;
  LUT3 id02064 (
    .ADR0(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[20].u_compressor42_cell.x2 ),
    .O(id04559)
  );

  defparam id02065.INIT = 8'hB2;
  LUT3 id02065 (
    .ADR0(id04144),
    .ADR1(id04149),
    .ADR2(id04150),
    .O(id04567)
  );

  defparam id02066.INIT = 8'h69;
  LUT3 id02066 (
    .ADR0(id04560),
    .ADR1(id04557),
    .ADR2(id04558),
    .O(\net_Buf-pad-result[22] )
  );

  defparam id02067.INIT = 16'hBF00;
  LUT4 id02067 (
    .ADR0(id04160),
    .ADR1(id04165),
    .ADR2(id04583),
    .ADR3(id04611),
    .O(id04560)
  );

  defparam id02068.INIT = 8'h17;
  LUT3 id02068 (
    .ADR0(id04578),
    .ADR1(id04584),
    .ADR2(id04581),
    .O(id04611)
  );

  defparam id02069.INIT = 4'h4;
  LUT2 id02069 (
    .ADR0(id04582),
    .ADR1(id04571),
    .O(id04557)
  );

  defparam id02070.INIT = 4'h9;
  LUT2 id02070 (
    .ADR0(id04612),
    .ADR1(id04609),
    .O(id04558)
  );

  defparam id02071.INIT = 8'hB2;
  LUT3 id02071 (
    .ADR0(id04572),
    .ADR1(id04570),
    .ADR2(id04569),
    .O(id04612)
  );

  defparam id02072.INIT = 4'h9;
  LUT2 id02072 (
    .ADR0(id04610),
    .ADR1(id04615),
    .O(id04609)
  );

  defparam id02073.INIT = 16'h9669;
  LUT4 id02073 (
    .ADR0(id04616),
    .ADR1(id04613),
    .ADR2(id04614),
    .ADR3(id04603),
    .O(id04610)
  );

  defparam id02074.INIT = 8'hC5;
  LUT3 id02074 (
    .ADR0(id04555),
    .ADR1(id04567),
    .ADR2(id04562),
    .O(id04616)
  );

  defparam id02075.INIT = 4'h9;
  LUT2 id02075 (
    .ADR0(id04604),
    .ADR1(id04601),
    .O(id04613)
  );

  defparam id02076.INIT = 16'h6996;
  LUT4 id02076 (
    .ADR0(id04602),
    .ADR1(id04607),
    .ADR2(id04608),
    .ADR3(id04605),
    .O(id04604)
  );

  defparam id02077.INIT = 8'h35;
  LUT3 id02077 (
    .ADR0(id04553),
    .ADR1(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x0 ),
    .ADR2(id04556),
    .O(id04602)
  );

  defparam id02078.INIT = 4'h9;
  LUT2 id02078 (
    .ADR0(id04606),
    .ADR1(id04595),
    .O(id04607)
  );

  defparam id02079.INIT = 16'h9669;
  LUT4 id02079 (
    .ADR0(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04606)
  );

  defparam id02080.INIT = 8'hE8;
  LUT3 id02080 (
    .ADR0(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04595)
  );

  defparam id02081.INIT = 16'h7117;
  LUT4 id02081 (
    .ADR0(id04559),
    .ADR1(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x0 ),
    .ADR2(id04554),
    .ADR3(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x3 ),
    .O(id04608)
  );

  defparam id02082.INIT = 16'h6996;
  LUT4 id02082 (
    .ADR0(id04596),
    .ADR1(id04593),
    .ADR2(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x3 ),
    .O(id04605)
  );

  defparam id02083.INIT = 4'h6;
  LUT2 id02083 (
    .ADR0(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x2 ),
    .O(id04596)
  );

  defparam id02084.INIT = 8'hE8;
  LUT3 id02084 (
    .ADR0(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[21].u_compressor42_cell.x2 ),
    .O(id04593)
  );

  defparam id02085.INIT = 8'hB2;
  LUT3 id02085 (
    .ADR0(id04568),
    .ADR1(id04565),
    .ADR2(id04566),
    .O(id04601)
  );

  defparam id02086.INIT = 4'h4;
  LUT2 id02086 (
    .ADR0(id04574),
    .ADR1(id04563),
    .O(id04614)
  );

  defparam id02087.INIT = 8'h69;
  LUT3 id02087 (
    .ADR0(id04594),
    .ADR1(id04599),
    .ADR2(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .O(id04603)
  );

  defparam id02088.INIT = 8'h35;
  LUT3 id02088 (
    .ADR0(id04561),
    .ADR1(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x0 ),
    .ADR2(id04564),
    .O(id04594)
  );

  defparam id02089.INIT = 4'h9;
  LUT2 id02089 (
    .ADR0(id04600),
    .ADR1(id04597),
    .O(id04599)
  );

  defparam id02090.INIT = 16'h9669;
  LUT4 id02090 (
    .ADR0(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04600)
  );

  defparam id02091.INIT = 8'hE8;
  LUT3 id02091 (
    .ADR0(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x1 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_2.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04597)
  );

  defparam id02092.INIT = 8'h2B;
  LUT3 id02092 (
    .ADR0(id04575),
    .ADR1(id04576),
    .ADR2(id04573),
    .O(id04615)
  );

  defparam id02093.INIT = 16'h2BD4;
  LUT4 id02093 (
    .ADR0(id04560),
    .ADR1(id04557),
    .ADR2(id04558),
    .ADR3(id04598),
    .O(\net_Buf-pad-result[23] )
  );

  defparam id02094.INIT = 4'h6;
  LUT2 id02094 (
    .ADR0(id04587),
    .ADR1(id04588),
    .O(id04598)
  );

  defparam id02095.INIT = 4'h4;
  LUT2 id02095 (
    .ADR0(id04612),
    .ADR1(id04609),
    .O(id04587)
  );

  defparam id02096.INIT = 4'h9;
  LUT2 id02096 (
    .ADR0(id04585),
    .ADR1(id04586),
    .O(id04588)
  );

  defparam id02097.INIT = 8'hC5;
  LUT3 id02097 (
    .ADR0(id04613),
    .ADR1(id04615),
    .ADR2(id04610),
    .O(id04585)
  );

  defparam id02098.INIT = 4'h6;
  LUT2 id02098 (
    .ADR0(id04591),
    .ADR1(id04592),
    .O(id04586)
  );

  defparam id02099.INIT = 16'h1EE1;
  LUT4 id02099 (
    .ADR0(id04589),
    .ADR1(id04590),
    .ADR2(id04515),
    .ADR3(id04516),
    .O(id04591)
  );

  defparam id02100.INIT = 16'h9000;
  LUT4 id02100 (
    .ADR0(id04594),
    .ADR1(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR2(id04599),
    .ADR3(id04513),
    .O(id04589)
  );

  defparam id02101.INIT = 8'h69;
  LUT3 id02101 (
    .ADR0(id04514),
    .ADR1(id04519),
    .ADR2(GND_NET),
    .O(id04513)
  );

  defparam id02102.INIT = 8'h35;
  LUT3 id02102 (
    .ADR0(id04597),
    .ADR1(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x0 ),
    .ADR2(id04600),
    .O(id04514)
  );

  defparam id02103.INIT = 16'h6996;
  LUT4 id02103 (
    .ADR0(id04520),
    .ADR1(id04517),
    .ADR2(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x3 ),
    .O(id04519)
  );

  defparam id02104.INIT = 4'h6;
  LUT2 id02104 (
    .ADR0(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04520)
  );

  defparam id02105.INIT = 8'hE8;
  LUT3 id02105 (
    .ADR0(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04517)
  );

  defparam id02106.INIT = 16'h304D;
  LUT4 id02106 (
    .ADR0(id04599),
    .ADR1(id04594),
    .ADR2(\DECODE_GEN[11].u_booth_enc.partial_reverse ),
    .ADR3(id04513),
    .O(id04590)
  );

  defparam id02107.INIT = 8'hC5;
  LUT3 id02107 (
    .ADR0(id04605),
    .ADR1(id04601),
    .ADR2(id04604),
    .O(id04515)
  );

  defparam id02108.INIT = 4'h6;
  LUT2 id02108 (
    .ADR0(id04518),
    .ADR1(id04507),
    .O(id04516)
  );

  defparam id02109.INIT = 16'h6996;
  LUT4 id02109 (
    .ADR0(id04508),
    .ADR1(id04505),
    .ADR2(id04506),
    .ADR3(id04511),
    .O(id04518)
  );

  defparam id02110.INIT = 8'h35;
  LUT3 id02110 (
    .ADR0(id04595),
    .ADR1(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x0 ),
    .ADR2(id04606),
    .O(id04508)
  );

  defparam id02111.INIT = 4'h9;
  LUT2 id02111 (
    .ADR0(id04512),
    .ADR1(id04509),
    .O(id04505)
  );

  defparam id02112.INIT = 16'h9669;
  LUT4 id02112 (
    .ADR0(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04512)
  );

  defparam id02113.INIT = 8'hE8;
  LUT3 id02113 (
    .ADR0(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04509)
  );

  defparam id02114.INIT = 16'h7117;
  LUT4 id02114 (
    .ADR0(id04593),
    .ADR1(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x0 ),
    .ADR2(id04596),
    .ADR3(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x3 ),
    .O(id04506)
  );

  defparam id02115.INIT = 16'h6996;
  LUT4 id02115 (
    .ADR0(id04510),
    .ADR1(id04499),
    .ADR2(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x3 ),
    .O(id04511)
  );

  defparam id02116.INIT = 4'h6;
  LUT2 id02116 (
    .ADR0(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x2 ),
    .O(id04510)
  );

  defparam id02117.INIT = 8'hE8;
  LUT3 id02117 (
    .ADR0(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[22].u_compressor42_cell.x2 ),
    .O(id04499)
  );

  defparam id02118.INIT = 8'h71;
  LUT3 id02118 (
    .ADR0(id04602),
    .ADR1(id04608),
    .ADR2(id04607),
    .O(id04507)
  );

  defparam id02119.INIT = 8'h2B;
  LUT3 id02119 (
    .ADR0(id04616),
    .ADR1(id04614),
    .ADR2(id04603),
    .O(id04592)
  );

  defparam id02120.INIT = 16'hE11E;
  LUT4 id02120 (
    .ADR0(id04500),
    .ADR1(id04497),
    .ADR2(id04498),
    .ADR3(id04503),
    .O(\net_Buf-pad-result[24] )
  );

  defparam id02121.INIT = 16'hD400;
  LUT4 id02121 (
    .ADR0(id04560),
    .ADR1(id04557),
    .ADR2(id04558),
    .ADR3(id04598),
    .O(id04500)
  );

  defparam id02122.INIT = 4'h8;
  LUT2 id02122 (
    .ADR0(id04587),
    .ADR1(id04588),
    .O(id04497)
  );

  defparam id02123.INIT = 4'h4;
  LUT2 id02123 (
    .ADR0(id04585),
    .ADR1(id04586),
    .O(id04498)
  );

  defparam id02124.INIT = 4'h9;
  LUT2 id02124 (
    .ADR0(id04504),
    .ADR1(id04501),
    .O(id04503)
  );

  defparam id02125.INIT = 8'h3A;
  LUT3 id02125 (
    .ADR0(id04592),
    .ADR1(id04516),
    .ADR2(id04591),
    .O(id04504)
  );

  defparam id02126.INIT = 4'h6;
  LUT2 id02126 (
    .ADR0(id04502),
    .ADR1(id04491),
    .O(id04501)
  );

  defparam id02127.INIT = 16'h6996;
  LUT4 id02127 (
    .ADR0(id04492),
    .ADR1(id04489),
    .ADR2(id04490),
    .ADR3(id04495),
    .O(id04502)
  );

  defparam id02128.INIT = 16'h1771;
  LUT4 id02128 (
    .ADR0(id04519),
    .ADR1(id04590),
    .ADR2(id04514),
    .ADR3(GND_NET),
    .O(id04492)
  );

  defparam id02129.INIT = 8'h96;
  LUT3 id02129 (
    .ADR0(id04496),
    .ADR1(id04493),
    .ADR2(id04494),
    .O(id04489)
  );

  defparam id02130.INIT = 4'h4;
  LUT2 id02130 (
    .ADR0(id04514),
    .ADR1(GND_NET),
    .O(id04496)
  );

  defparam id02131.INIT = 8'h69;
  LUT3 id02131 (
    .ADR0(id04547),
    .ADR1(\u_compressor42_l0_3.CELLS[2].u_compressor42_cell.x0 ),
    .ADR2(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .O(id04493)
  );

  defparam id02132.INIT = 16'h7117;
  LUT4 id02132 (
    .ADR0(id04517),
    .ADR1(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x0 ),
    .ADR2(id04520),
    .ADR3(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x3 ),
    .O(id04547)
  );

  defparam id02133.INIT = 16'h6996;
  LUT4 id02133 (
    .ADR0(id04548),
    .ADR1(id04545),
    .ADR2(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x3 ),
    .O(id04494)
  );

  defparam id02134.INIT = 4'h6;
  LUT2 id02134 (
    .ADR0(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04548)
  );

  defparam id02135.INIT = 8'hE8;
  LUT3 id02135 (
    .ADR0(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04545)
  );

  defparam id02136.INIT = 8'h35;
  LUT3 id02136 (
    .ADR0(id04511),
    .ADR1(id04507),
    .ADR2(id04518),
    .O(id04490)
  );

  defparam id02137.INIT = 4'h9;
  LUT2 id02137 (
    .ADR0(id04546),
    .ADR1(id04551),
    .O(id04495)
  );

  defparam id02138.INIT = 16'h6996;
  LUT4 id02138 (
    .ADR0(id04552),
    .ADR1(id04549),
    .ADR2(id04550),
    .ADR3(id04539),
    .O(id04546)
  );

  defparam id02139.INIT = 8'h35;
  LUT3 id02139 (
    .ADR0(id04509),
    .ADR1(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x0 ),
    .ADR2(id04512),
    .O(id04552)
  );

  defparam id02140.INIT = 4'h9;
  LUT2 id02140 (
    .ADR0(id04540),
    .ADR1(id04537),
    .O(id04549)
  );

  defparam id02141.INIT = 16'h9669;
  LUT4 id02141 (
    .ADR0(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x2 ),
    .O(id04540)
  );

  defparam id02142.INIT = 8'hE8;
  LUT3 id02142 (
    .ADR0(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04537)
  );

  defparam id02143.INIT = 16'h7117;
  LUT4 id02143 (
    .ADR0(id04499),
    .ADR1(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x0 ),
    .ADR2(id04510),
    .ADR3(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x3 ),
    .O(id04550)
  );

  defparam id02144.INIT = 16'h6996;
  LUT4 id02144 (
    .ADR0(id04538),
    .ADR1(id04543),
    .ADR2(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x3 ),
    .O(id04539)
  );

  defparam id02145.INIT = 4'h6;
  LUT2 id02145 (
    .ADR0(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x2 ),
    .O(id04538)
  );

  defparam id02146.INIT = 8'hE8;
  LUT3 id02146 (
    .ADR0(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[23].u_compressor42_cell.x2 ),
    .O(id04543)
  );

  defparam id02147.INIT = 8'hB2;
  LUT3 id02147 (
    .ADR0(id04508),
    .ADR1(id04505),
    .ADR2(id04506),
    .O(id04551)
  );

  defparam id02148.INIT = 8'h0D;
  LUT3 id02148 (
    .ADR0(id04515),
    .ADR1(id04589),
    .ADR2(id04590),
    .O(id04491)
  );

  defparam id02149.INIT = 8'h69;
  LUT3 id02149 (
    .ADR0(id04544),
    .ADR1(id04541),
    .ADR2(id04542),
    .O(\net_Buf-pad-result[25] )
  );

  defparam id02150.INIT = 16'h1117;
  LUT4 id02150 (
    .ADR0(id04498),
    .ADR1(id04503),
    .ADR2(id04500),
    .ADR3(id04497),
    .O(id04544)
  );

  defparam id02151.INIT = 4'h4;
  LUT2 id02151 (
    .ADR0(id04504),
    .ADR1(id04501),
    .O(id04541)
  );

  defparam id02152.INIT = 4'h9;
  LUT2 id02152 (
    .ADR0(id04531),
    .ADR1(id04532),
    .O(id04542)
  );

  defparam id02153.INIT = 8'h35;
  LUT3 id02153 (
    .ADR0(id04495),
    .ADR1(id04491),
    .ADR2(id04502),
    .O(id04531)
  );

  defparam id02154.INIT = 4'h9;
  LUT2 id02154 (
    .ADR0(id04529),
    .ADR1(id04530),
    .O(id04532)
  );

  defparam id02155.INIT = 16'h6996;
  LUT4 id02155 (
    .ADR0(id04535),
    .ADR1(id04536),
    .ADR2(id04533),
    .ADR3(id04534),
    .O(id04529)
  );

  defparam id02156.INIT = 8'h17;
  LUT3 id02156 (
    .ADR0(id04496),
    .ADR1(id04493),
    .ADR2(id04494),
    .O(id04535)
  );

  defparam id02157.INIT = 16'h9669;
  LUT4 id02157 (
    .ADR0(id04523),
    .ADR1(id04524),
    .ADR2(id04521),
    .ADR3(id04522),
    .O(id04536)
  );

  defparam id02158.INIT = 8'h14;
  LUT3 id02158 (
    .ADR0(id04547),
    .ADR1(\u_compressor42_l0_3.CELLS[2].u_compressor42_cell.x0 ),
    .ADR2(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .O(id04523)
  );

  defparam id02159.INIT = 16'h6996;
  LUT4 id02159 (
    .ADR0(id04527),
    .ADR1(id04528),
    .ADR2(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x3 ),
    .O(id04524)
  );

  defparam id02160.INIT = 4'h6;
  LUT2 id02160 (
    .ADR0(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x2 ),
    .O(id04527)
  );

  defparam id02161.INIT = 8'hE8;
  LUT3 id02161 (
    .ADR0(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04528)
  );

  defparam id02162.INIT = 16'h7117;
  LUT4 id02162 (
    .ADR0(id04545),
    .ADR1(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x0 ),
    .ADR2(id04548),
    .ADR3(\u_compressor42_l0_2.CELLS[10].u_compressor42_cell.x3 ),
    .O(id04521)
  );

  defparam id02163.INIT = 8'h96;
  LUT3 id02163 (
    .ADR0(id04525),
    .ADR1(\u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .O(id04522)
  );

  defparam id02164.INIT = 4'h8;
  LUT2 id02164 (
    .ADR0(\u_compressor42_l0_3.CELLS[2].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[12].u_booth_enc.partial_reverse ),
    .O(id04525)
  );

  defparam id02165.INIT = 8'hC5;
  LUT3 id02165 (
    .ADR0(id04539),
    .ADR1(id04551),
    .ADR2(id04546),
    .O(id04533)
  );

  defparam id02166.INIT = 4'h6;
  LUT2 id02166 (
    .ADR0(id04526),
    .ADR1(id04707),
    .O(id04534)
  );

  defparam id02167.INIT = 16'h9669;
  LUT4 id02167 (
    .ADR0(id04708),
    .ADR1(id04705),
    .ADR2(id04706),
    .ADR3(id04711),
    .O(id04526)
  );

  defparam id02168.INIT = 8'h35;
  LUT3 id02168 (
    .ADR0(id04537),
    .ADR1(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x0 ),
    .ADR2(id04540),
    .O(id04708)
  );

  defparam id02169.INIT = 4'h9;
  LUT2 id02169 (
    .ADR0(id04712),
    .ADR1(id04709),
    .O(id04705)
  );

  defparam id02170.INIT = 16'h9669;
  LUT4 id02170 (
    .ADR0(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x2 ),
    .O(id04712)
  );

  defparam id02171.INIT = 8'hE8;
  LUT3 id02171 (
    .ADR0(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[18].u_compressor42_cell.x2 ),
    .O(id04709)
  );

  defparam id02172.INIT = 16'h7117;
  LUT4 id02172 (
    .ADR0(id04543),
    .ADR1(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x0 ),
    .ADR2(id04538),
    .ADR3(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x3 ),
    .O(id04706)
  );

  defparam id02173.INIT = 16'h6996;
  LUT4 id02173 (
    .ADR0(id04710),
    .ADR1(id04699),
    .ADR2(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x3 ),
    .O(id04711)
  );

  defparam id02174.INIT = 4'h6;
  LUT2 id02174 (
    .ADR0(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x2 ),
    .O(id04710)
  );

  defparam id02175.INIT = 8'hE8;
  LUT3 id02175 (
    .ADR0(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[24].u_compressor42_cell.x2 ),
    .O(id04699)
  );

  defparam id02176.INIT = 8'hB2;
  LUT3 id02176 (
    .ADR0(id04552),
    .ADR1(id04549),
    .ADR2(id04550),
    .O(id04707)
  );

  defparam id02177.INIT = 8'hB2;
  LUT3 id02177 (
    .ADR0(id04492),
    .ADR1(id04489),
    .ADR2(id04490),
    .O(id04530)
  );

  defparam id02178.INIT = 16'h2BD4;
  LUT4 id02178 (
    .ADR0(id04544),
    .ADR1(id04541),
    .ADR2(id04542),
    .ADR3(id04700),
    .O(\net_Buf-pad-result[26] )
  );

  defparam id02179.INIT = 4'h6;
  LUT2 id02179 (
    .ADR0(id04697),
    .ADR1(id04698),
    .O(id04700)
  );

  defparam id02180.INIT = 4'h4;
  LUT2 id02180 (
    .ADR0(id04531),
    .ADR1(id04532),
    .O(id04697)
  );

  defparam id02181.INIT = 4'h9;
  LUT2 id02181 (
    .ADR0(id04703),
    .ADR1(id04704),
    .O(id04698)
  );

  defparam id02182.INIT = 8'hC5;
  LUT3 id02182 (
    .ADR0(id04534),
    .ADR1(id04530),
    .ADR2(id04529),
    .O(id04703)
  );

  defparam id02183.INIT = 4'h9;
  LUT2 id02183 (
    .ADR0(id04701),
    .ADR1(id04702),
    .O(id04704)
  );

  defparam id02184.INIT = 16'h9669;
  LUT4 id02184 (
    .ADR0(id04691),
    .ADR1(id04692),
    .ADR2(id04689),
    .ADR3(id04690),
    .O(id04701)
  );

  defparam id02185.INIT = 16'h1771;
  LUT4 id02185 (
    .ADR0(id04523),
    .ADR1(id04524),
    .ADR2(id04521),
    .ADR3(id04522),
    .O(id04691)
  );

  defparam id02186.INIT = 8'h69;
  LUT3 id02186 (
    .ADR0(id04695),
    .ADR1(id04696),
    .ADR2(id04693),
    .O(id04692)
  );

  defparam id02187.INIT = 16'h8778;
  LUT4 id02187 (
    .ADR0(\u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(id04694),
    .ADR3(id04683),
    .O(id04695)
  );

  defparam id02188.INIT = 16'h6996;
  LUT4 id02188 (
    .ADR0(id04684),
    .ADR1(id04681),
    .ADR2(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x3 ),
    .O(id04694)
  );

  defparam id02189.INIT = 4'h6;
  LUT2 id02189 (
    .ADR0(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x2 ),
    .O(id04684)
  );

  defparam id02190.INIT = 8'hE8;
  LUT3 id02190 (
    .ADR0(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x2 ),
    .O(id04681)
  );

  defparam id02191.INIT = 8'h96;
  LUT3 id02191 (
    .ADR0(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 ),
    .O(id04683)
  );

  defparam id02192.INIT = 16'hB22B;
  LUT4 id02192 (
    .ADR0(id04521),
    .ADR1(id04525),
    .ADR2(\u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04696)
  );

  defparam id02193.INIT = 16'h7117;
  LUT4 id02193 (
    .ADR0(id04528),
    .ADR1(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x0 ),
    .ADR2(id04527),
    .ADR3(\u_compressor42_l0_2.CELLS[11].u_compressor42_cell.x3 ),
    .O(id04693)
  );

  defparam id02194.INIT = 8'h3A;
  LUT3 id02194 (
    .ADR0(id04707),
    .ADR1(id04711),
    .ADR2(id04526),
    .O(id04689)
  );

  defparam id02195.INIT = 4'h6;
  LUT2 id02195 (
    .ADR0(id04682),
    .ADR1(id04687),
    .O(id04690)
  );

  defparam id02196.INIT = 16'h6996;
  LUT4 id02196 (
    .ADR0(id04688),
    .ADR1(id04685),
    .ADR2(id04686),
    .ADR3(id04739),
    .O(id04682)
  );

  defparam id02197.INIT = 8'h35;
  LUT3 id02197 (
    .ADR0(id04709),
    .ADR1(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x0 ),
    .ADR2(id04712),
    .O(id04688)
  );

  defparam id02198.INIT = 4'h9;
  LUT2 id02198 (
    .ADR0(id04740),
    .ADR1(id04737),
    .O(id04685)
  );

  defparam id02199.INIT = 16'h9669;
  LUT4 id02199 (
    .ADR0(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x2 ),
    .O(id04740)
  );

  defparam id02200.INIT = 8'hE8;
  LUT3 id02200 (
    .ADR0(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[19].u_compressor42_cell.x2 ),
    .O(id04737)
  );

  defparam id02201.INIT = 16'h7117;
  LUT4 id02201 (
    .ADR0(id04699),
    .ADR1(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x0 ),
    .ADR2(id04710),
    .ADR3(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x3 ),
    .O(id04686)
  );

  defparam id02202.INIT = 16'h6996;
  LUT4 id02202 (
    .ADR0(id04738),
    .ADR1(id04743),
    .ADR2(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x3 ),
    .O(id04739)
  );

  defparam id02203.INIT = 4'h6;
  LUT2 id02203 (
    .ADR0(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x2 ),
    .O(id04738)
  );

  defparam id02204.INIT = 8'hE8;
  LUT3 id02204 (
    .ADR0(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[25].u_compressor42_cell.x2 ),
    .O(id04743)
  );

  defparam id02205.INIT = 8'h71;
  LUT3 id02205 (
    .ADR0(id04708),
    .ADR1(id04706),
    .ADR2(id04705),
    .O(id04687)
  );

  defparam id02206.INIT = 8'hB2;
  LUT3 id02206 (
    .ADR0(id04535),
    .ADR1(id04536),
    .ADR2(id04533),
    .O(id04702)
  );

  defparam id02207.INIT = 8'h1E;
  LUT3 id02207 (
    .ADR0(id04744),
    .ADR1(id04741),
    .ADR2(id04742),
    .O(\net_Buf-pad-result[27] )
  );

  defparam id02208.INIT = 16'hD400;
  LUT4 id02208 (
    .ADR0(id04544),
    .ADR1(id04541),
    .ADR2(id04542),
    .ADR3(id04700),
    .O(id04744)
  );

  defparam id02209.INIT = 4'h8;
  LUT2 id02209 (
    .ADR0(id04697),
    .ADR1(id04698),
    .O(id04741)
  );

  defparam id02210.INIT = 4'h6;
  LUT2 id02210 (
    .ADR0(id04731),
    .ADR1(id04732),
    .O(id04742)
  );

  defparam id02211.INIT = 4'h4;
  LUT2 id02211 (
    .ADR0(id04703),
    .ADR1(id04704),
    .O(id04731)
  );

  defparam id02212.INIT = 4'h9;
  LUT2 id02212 (
    .ADR0(id04729),
    .ADR1(id04730),
    .O(id04732)
  );

  defparam id02213.INIT = 8'hC5;
  LUT3 id02213 (
    .ADR0(id04690),
    .ADR1(id04702),
    .ADR2(id04701),
    .O(id04729)
  );

  defparam id02214.INIT = 4'h9;
  LUT2 id02214 (
    .ADR0(id04735),
    .ADR1(id04736),
    .O(id04730)
  );

  defparam id02215.INIT = 16'h9669;
  LUT4 id02215 (
    .ADR0(id04733),
    .ADR1(id04734),
    .ADR2(id04723),
    .ADR3(id04724),
    .O(id04735)
  );

  defparam id02216.INIT = 16'h5CC5;
  LUT4 id02216 (
    .ADR0(id04696),
    .ADR1(id04694),
    .ADR2(id04695),
    .ADR3(id04693),
    .O(id04733)
  );

  defparam id02217.INIT = 4'h9;
  LUT2 id02217 (
    .ADR0(id04721),
    .ADR1(id04722),
    .O(id04734)
  );

  defparam id02218.INIT = 16'hE11E;
  LUT4 id02218 (
    .ADR0(id04727),
    .ADR1(id04728),
    .ADR2(id04725),
    .ADR3(id04726),
    .O(id04721)
  );

  defparam id02219.INIT = 16'h6000;
  LUT4 id02219 (
    .ADR0(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 ),
    .ADR2(id04715),
    .ADR3(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x0 ),
    .O(id04727)
  );

  defparam id02220.INIT = 8'h96;
  LUT3 id02220 (
    .ADR0(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x0 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 ),
    .O(id04715)
  );

  defparam id02221.INIT = 16'hC017;
  LUT4 id02221 (
    .ADR0(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x0 ),
    .ADR1(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 ),
    .ADR3(id04715),
    .O(id04728)
  );

  defparam id02222.INIT = 16'h7117;
  LUT4 id02222 (
    .ADR0(id04681),
    .ADR1(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x0 ),
    .ADR2(id04684),
    .ADR3(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x3 ),
    .O(id04725)
  );

  defparam id02223.INIT = 16'h6996;
  LUT4 id02223 (
    .ADR0(id04716),
    .ADR1(id04713),
    .ADR2(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x3 ),
    .O(id04726)
  );

  defparam id02224.INIT = 4'h6;
  LUT2 id02224 (
    .ADR0(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04716)
  );

  defparam id02225.INIT = 8'hE8;
  LUT3 id02225 (
    .ADR0(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[12].u_compressor42_cell.x2 ),
    .O(id04713)
  );

  defparam id02226.INIT = 16'h2BBB;
  LUT4 id02226 (
    .ADR0(id04693),
    .ADR1(id04683),
    .ADR2(\u_compressor42_l0_3.CELLS[3].u_compressor42_cell.x0 ),
    .ADR3(GND_NET),
    .O(id04722)
  );

  defparam id02227.INIT = 8'h35;
  LUT3 id02227 (
    .ADR0(id04739),
    .ADR1(id04687),
    .ADR2(id04682),
    .O(id04723)
  );

  defparam id02228.INIT = 4'h6;
  LUT2 id02228 (
    .ADR0(id04714),
    .ADR1(id04719),
    .O(id04724)
  );

  defparam id02229.INIT = 16'h6996;
  LUT4 id02229 (
    .ADR0(id04720),
    .ADR1(id04717),
    .ADR2(id04718),
    .ADR3(id04643),
    .O(id04714)
  );

  defparam id02230.INIT = 8'h35;
  LUT3 id02230 (
    .ADR0(id04737),
    .ADR1(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x0 ),
    .ADR2(id04740),
    .O(id04720)
  );

  defparam id02231.INIT = 4'h9;
  LUT2 id02231 (
    .ADR0(id04644),
    .ADR1(id04641),
    .O(id04717)
  );

  defparam id02232.INIT = 16'h9669;
  LUT4 id02232 (
    .ADR0(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x2 ),
    .O(id04644)
  );

  defparam id02233.INIT = 8'hE8;
  LUT3 id02233 (
    .ADR0(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[20].u_compressor42_cell.x2 ),
    .O(id04641)
  );

  defparam id02234.INIT = 16'h7117;
  LUT4 id02234 (
    .ADR0(id04743),
    .ADR1(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x0 ),
    .ADR2(id04738),
    .ADR3(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x3 ),
    .O(id04718)
  );

  defparam id02235.INIT = 16'h6996;
  LUT4 id02235 (
    .ADR0(id04642),
    .ADR1(id04647),
    .ADR2(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x3 ),
    .O(id04643)
  );

  defparam id02236.INIT = 4'h6;
  LUT2 id02236 (
    .ADR0(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x2 ),
    .O(id04642)
  );

  defparam id02237.INIT = 8'hE8;
  LUT3 id02237 (
    .ADR0(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[26].u_compressor42_cell.x2 ),
    .O(id04647)
  );

  defparam id02238.INIT = 8'h71;
  LUT3 id02238 (
    .ADR0(id04688),
    .ADR1(id04686),
    .ADR2(id04685),
    .O(id04719)
  );

  defparam id02239.INIT = 8'hE8;
  LUT3 id02239 (
    .ADR0(id04691),
    .ADR1(id04692),
    .ADR2(id04689),
    .O(id04736)
  );

  defparam id02240.INIT = 16'h07F8;
  LUT4 id02240 (
    .ADR0(id04744),
    .ADR1(id04742),
    .ADR2(id04648),
    .ADR3(id04645),
    .O(\net_Buf-pad-result[28] )
  );

  defparam id02241.INIT = 8'hE0;
  LUT3 id02241 (
    .ADR0(id04731),
    .ADR1(id04741),
    .ADR2(id04732),
    .O(id04648)
  );

  defparam id02242.INIT = 4'h6;
  LUT2 id02242 (
    .ADR0(id04646),
    .ADR1(id04635),
    .O(id04645)
  );

  defparam id02243.INIT = 4'h4;
  LUT2 id02243 (
    .ADR0(id04729),
    .ADR1(id04730),
    .O(id04646)
  );

  defparam id02244.INIT = 4'h9;
  LUT2 id02244 (
    .ADR0(id04636),
    .ADR1(id04633),
    .O(id04635)
  );

  defparam id02245.INIT = 8'hC5;
  LUT3 id02245 (
    .ADR0(id04724),
    .ADR1(id04736),
    .ADR2(id04735),
    .O(id04636)
  );

  defparam id02246.INIT = 4'h9;
  LUT2 id02246 (
    .ADR0(id04634),
    .ADR1(id04639),
    .O(id04633)
  );

  defparam id02247.INIT = 16'h9669;
  LUT4 id02247 (
    .ADR0(id04640),
    .ADR1(id04637),
    .ADR2(id04638),
    .ADR3(id04627),
    .O(id04634)
  );

  defparam id02248.INIT = 8'hC5;
  LUT3 id02248 (
    .ADR0(id04726),
    .ADR1(id04722),
    .ADR2(id04721),
    .O(id04640)
  );

  defparam id02249.INIT = 4'h6;
  LUT2 id02249 (
    .ADR0(id04628),
    .ADR1(id04625),
    .O(id04637)
  );

  defparam id02250.INIT = 16'h6996;
  LUT4 id02250 (
    .ADR0(id04626),
    .ADR1(id04631),
    .ADR2(id04632),
    .ADR3(id04629),
    .O(id04628)
  );

  defparam id02251.INIT = 16'h7117;
  LUT4 id02251 (
    .ADR0(id04630),
    .ADR1(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x0 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 ),
    .O(id04626)
  );

  defparam id02252.INIT = 4'h8;
  LUT2 id02252 (
    .ADR0(\DECODE_GEN[13].u_booth_enc.partial_reverse ),
    .ADR1(\u_compressor42_l0_3.CELLS[4].u_compressor42_cell.x1 ),
    .O(id04630)
  );

  defparam id02253.INIT = 8'h87;
  LUT3 id02253 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(id04619),
    .O(id04631)
  );

  defparam id02254.INIT = 16'h9669;
  LUT4 id02254 (
    .ADR0(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x1 ),
    .ADR2(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR3(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04619)
  );

  defparam id02255.INIT = 16'h7117;
  LUT4 id02255 (
    .ADR0(id04713),
    .ADR1(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x0 ),
    .ADR2(id04716),
    .ADR3(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x3 ),
    .O(id04632)
  );

  defparam id02256.INIT = 16'h6996;
  LUT4 id02256 (
    .ADR0(id04620),
    .ADR1(id04617),
    .ADR2(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x3 ),
    .O(id04629)
  );

  defparam id02257.INIT = 4'h6;
  LUT2 id02257 (
    .ADR0(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04620)
  );

  defparam id02258.INIT = 8'hE8;
  LUT3 id02258 (
    .ADR0(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[13].u_compressor42_cell.x2 ),
    .O(id04617)
  );

  defparam id02259.INIT = 8'h0D;
  LUT3 id02259 (
    .ADR0(id04725),
    .ADR1(id04727),
    .ADR2(id04728),
    .O(id04625)
  );

  defparam id02260.INIT = 8'h35;
  LUT3 id02260 (
    .ADR0(id04643),
    .ADR1(id04719),
    .ADR2(id04714),
    .O(id04638)
  );

  defparam id02261.INIT = 4'h9;
  LUT2 id02261 (
    .ADR0(id04618),
    .ADR1(id04623),
    .O(id04627)
  );

  defparam id02262.INIT = 16'h6996;
  LUT4 id02262 (
    .ADR0(id04624),
    .ADR1(id04621),
    .ADR2(id04622),
    .ADR3(id04675),
    .O(id04618)
  );

  defparam id02263.INIT = 8'h35;
  LUT3 id02263 (
    .ADR0(id04641),
    .ADR1(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x0 ),
    .ADR2(id04644),
    .O(id04624)
  );

  defparam id02264.INIT = 4'h9;
  LUT2 id02264 (
    .ADR0(id04676),
    .ADR1(id04673),
    .O(id04621)
  );

  defparam id02265.INIT = 16'h9669;
  LUT4 id02265 (
    .ADR0(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x2 ),
    .O(id04676)
  );

  defparam id02266.INIT = 8'hE8;
  LUT3 id02266 (
    .ADR0(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[21].u_compressor42_cell.x2 ),
    .O(id04673)
  );

  defparam id02267.INIT = 16'h7117;
  LUT4 id02267 (
    .ADR0(id04647),
    .ADR1(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x0 ),
    .ADR2(id04642),
    .ADR3(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x3 ),
    .O(id04622)
  );

  defparam id02268.INIT = 16'h6996;
  LUT4 id02268 (
    .ADR0(id04674),
    .ADR1(id04679),
    .ADR2(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x3 ),
    .O(id04675)
  );

  defparam id02269.INIT = 4'h6;
  LUT2 id02269 (
    .ADR0(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x2 ),
    .O(id04674)
  );

  defparam id02270.INIT = 8'hE8;
  LUT3 id02270 (
    .ADR0(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[27].u_compressor42_cell.x2 ),
    .O(id04679)
  );

  defparam id02271.INIT = 8'hB2;
  LUT3 id02271 (
    .ADR0(id04720),
    .ADR1(id04717),
    .ADR2(id04718),
    .O(id04623)
  );

  defparam id02272.INIT = 8'hB2;
  LUT3 id02272 (
    .ADR0(id04733),
    .ADR1(id04723),
    .ADR2(id04734),
    .O(id04639)
  );

  defparam id02273.INIT = 8'h1E;
  LUT3 id02273 (
    .ADR0(id04680),
    .ADR1(id04677),
    .ADR2(id04678),
    .O(\net_Buf-pad-result[29] )
  );

  defparam id02274.INIT = 16'hF800;
  LUT4 id02274 (
    .ADR0(id04744),
    .ADR1(id04742),
    .ADR2(id04648),
    .ADR3(id04645),
    .O(id04680)
  );

  defparam id02275.INIT = 4'h8;
  LUT2 id02275 (
    .ADR0(id04646),
    .ADR1(id04635),
    .O(id04677)
  );

  defparam id02276.INIT = 4'h6;
  LUT2 id02276 (
    .ADR0(id04667),
    .ADR1(id04668),
    .O(id04678)
  );

  defparam id02277.INIT = 4'h4;
  LUT2 id02277 (
    .ADR0(id04636),
    .ADR1(id04633),
    .O(id04667)
  );

  defparam id02278.INIT = 4'h9;
  LUT2 id02278 (
    .ADR0(id04665),
    .ADR1(id04666),
    .O(id04668)
  );

  defparam id02279.INIT = 8'h35;
  LUT3 id02279 (
    .ADR0(id04639),
    .ADR1(id04627),
    .ADR2(id04634),
    .O(id04665)
  );

  defparam id02280.INIT = 4'h6;
  LUT2 id02280 (
    .ADR0(id04671),
    .ADR1(id04672),
    .O(id04666)
  );

  defparam id02281.INIT = 16'h9669;
  LUT4 id02281 (
    .ADR0(id04669),
    .ADR1(id04670),
    .ADR2(id04659),
    .ADR3(id04660),
    .O(id04671)
  );

  defparam id02282.INIT = 8'h35;
  LUT3 id02282 (
    .ADR0(id04629),
    .ADR1(id04625),
    .ADR2(id04628),
    .O(id04669)
  );

  defparam id02283.INIT = 4'h6;
  LUT2 id02283 (
    .ADR0(id04657),
    .ADR1(id04658),
    .O(id04670)
  );

  defparam id02284.INIT = 16'h6996;
  LUT4 id02284 (
    .ADR0(id04663),
    .ADR1(id04664),
    .ADR2(id04661),
    .ADR3(id04662),
    .O(id04657)
  );

  defparam id02285.INIT = 16'h0F77;
  LUT4 id02285 (
    .ADR0(GND_NET),
    .ADR1(\u_compressor42_l0_3.CELLS[5].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x0 ),
    .ADR3(id04619),
    .O(id04663)
  );

  defparam id02286.INIT = 4'h9;
  LUT2 id02286 (
    .ADR0(id04651),
    .ADR1(id04652),
    .O(id04664)
  );

  defparam id02287.INIT = 16'h9669;
  LUT4 id02287 (
    .ADR0(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x1 ),
    .ADR2(GND_NET),
    .ADR3(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04651)
  );

  defparam id02288.INIT = 8'hE8;
  LUT3 id02288 (
    .ADR0(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x1 ),
    .ADR1(\DECODE_GEN[14].u_booth_enc.partial_reverse ),
    .ADR2(\u_compressor42_l0_3.CELLS[6].u_compressor42_cell.x2 ),
    .O(id04652)
  );

  defparam id02289.INIT = 16'h7117;
  LUT4 id02289 (
    .ADR0(id04617),
    .ADR1(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x0 ),
    .ADR2(id04620),
    .ADR3(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x3 ),
    .O(id04661)
  );

  defparam id02290.INIT = 16'h6996;
  LUT4 id02290 (
    .ADR0(id04649),
    .ADR1(id04650),
    .ADR2(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x3 ),
    .O(id04662)
  );

  defparam id02291.INIT = 4'h6;
  LUT2 id02291 (
    .ADR0(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04649)
  );

  defparam id02292.INIT = 8'hE8;
  LUT3 id02292 (
    .ADR0(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[14].u_compressor42_cell.x2 ),
    .O(id04650)
  );

  defparam id02293.INIT = 8'h71;
  LUT3 id02293 (
    .ADR0(id04626),
    .ADR1(id04632),
    .ADR2(id04631),
    .O(id04658)
  );

  defparam id02294.INIT = 8'hC5;
  LUT3 id02294 (
    .ADR0(id04675),
    .ADR1(id04623),
    .ADR2(id04618),
    .O(id04659)
  );

  defparam id02295.INIT = 4'h6;
  LUT2 id02295 (
    .ADR0(id04655),
    .ADR1(id04656),
    .O(id04660)
  );

  defparam id02296.INIT = 16'h9669;
  LUT4 id02296 (
    .ADR0(id04653),
    .ADR1(id04654),
    .ADR2(id04821),
    .ADR3(id04822),
    .O(id04655)
  );

  defparam id02297.INIT = 8'h35;
  LUT3 id02297 (
    .ADR0(id04673),
    .ADR1(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x0 ),
    .ADR2(id04676),
    .O(id04653)
  );

  defparam id02298.INIT = 4'h9;
  LUT2 id02298 (
    .ADR0(id04819),
    .ADR1(id04820),
    .O(id04654)
  );

  defparam id02299.INIT = 16'h9669;
  LUT4 id02299 (
    .ADR0(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x2 ),
    .O(id04819)
  );

  defparam id02300.INIT = 8'hE8;
  LUT3 id02300 (
    .ADR0(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[22].u_compressor42_cell.x2 ),
    .O(id04820)
  );

  defparam id02301.INIT = 16'h7117;
  LUT4 id02301 (
    .ADR0(id04679),
    .ADR1(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x0 ),
    .ADR2(id04674),
    .ADR3(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x3 ),
    .O(id04821)
  );

  defparam id02302.INIT = 16'h6996;
  LUT4 id02302 (
    .ADR0(id04825),
    .ADR1(id04826),
    .ADR2(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x3 ),
    .O(id04822)
  );

  defparam id02303.INIT = 4'h6;
  LUT2 id02303 (
    .ADR0(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x2 ),
    .O(id04825)
  );

  defparam id02304.INIT = 8'hE8;
  LUT3 id02304 (
    .ADR0(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[28].u_compressor42_cell.x2 ),
    .O(id04826)
  );

  defparam id02305.INIT = 8'hB2;
  LUT3 id02305 (
    .ADR0(id04624),
    .ADR1(id04621),
    .ADR2(id04622),
    .O(id04656)
  );

  defparam id02306.INIT = 8'hB2;
  LUT3 id02306 (
    .ADR0(id04640),
    .ADR1(id04637),
    .ADR2(id04638),
    .O(id04672)
  );

  defparam id02307.INIT = 4'h9;
  LUT2 id02307 (
    .ADR0(id04823),
    .ADR1(id04824),
    .O(\net_Buf-pad-result[30] )
  );

  defparam id02308.INIT = 16'h1117;
  LUT4 id02308 (
    .ADR0(id04667),
    .ADR1(id04668),
    .ADR2(id04680),
    .ADR3(id04677),
    .O(id04823)
  );

  defparam id02309.INIT = 4'h9;
  LUT2 id02309 (
    .ADR0(id04813),
    .ADR1(id04814),
    .O(id04824)
  );

  defparam id02310.INIT = 4'h4;
  LUT2 id02310 (
    .ADR0(id04665),
    .ADR1(id04666),
    .O(id04813)
  );

  defparam id02311.INIT = 8'h96;
  LUT3 id02311 (
    .ADR0(id04811),
    .ADR1(id04812),
    .ADR2(id03943),
    .O(id04814)
  );

  defparam id02312.INIT = 8'h3A;
  LUT3 id02312 (
    .ADR0(id04672),
    .ADR1(id04660),
    .ADR2(id04671),
    .O(id04811)
  );

  defparam id02313.INIT = 4'h9;
  LUT2 id02313 (
    .ADR0(id04817),
    .ADR1(id04818),
    .O(id04812)
  );

  defparam id02314.INIT = 16'h6996;
  LUT4 id02314 (
    .ADR0(id04815),
    .ADR1(id04816),
    .ADR2(id04805),
    .ADR3(id04806),
    .O(id04817)
  );

  defparam id02315.INIT = 8'h35;
  LUT3 id02315 (
    .ADR0(id04662),
    .ADR1(id04658),
    .ADR2(id04657),
    .O(id04815)
  );

  defparam id02316.INIT = 4'h6;
  LUT2 id02316 (
    .ADR0(id04803),
    .ADR1(id04804),
    .O(id04816)
  );

  defparam id02317.INIT = 16'h9669;
  LUT4 id02317 (
    .ADR0(id04809),
    .ADR1(id04810),
    .ADR2(id04807),
    .ADR3(id04808),
    .O(id04803)
  );

  defparam id02318.INIT = 8'h35;
  LUT3 id02318 (
    .ADR0(id04652),
    .ADR1(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x0 ),
    .ADR2(id04651),
    .O(id04809)
  );

  defparam id02319.INIT = 4'h9;
  LUT2 id02319 (
    .ADR0(id04797),
    .ADR1(id04798),
    .O(id04810)
  );

  defparam id02320.INIT = 16'h9669;
  LUT4 id02320 (
    .ADR0(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04797)
  );

  defparam id02321.INIT = 8'hE8;
  LUT3 id02321 (
    .ADR0(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x1 ),
    .ADR1(GND_NET),
    .ADR2(\u_compressor42_l0_3.CELLS[7].u_compressor42_cell.x2 ),
    .O(id04798)
  );

  defparam id02322.INIT = 16'h7117;
  LUT4 id02322 (
    .ADR0(id04650),
    .ADR1(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x0 ),
    .ADR2(id04649),
    .ADR3(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x3 ),
    .O(id04807)
  );

  defparam id02323.INIT = 16'h6996;
  LUT4 id02323 (
    .ADR0(id04795),
    .ADR1(id04796),
    .ADR2(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x3 ),
    .O(id04808)
  );

  defparam id02324.INIT = 4'h6;
  LUT2 id02324 (
    .ADR0(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04795)
  );

  defparam id02325.INIT = 8'hE8;
  LUT3 id02325 (
    .ADR0(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[15].u_compressor42_cell.x2 ),
    .O(id04796)
  );

  defparam id02326.INIT = 8'hB2;
  LUT3 id02326 (
    .ADR0(id04663),
    .ADR1(id04664),
    .ADR2(id04661),
    .O(id04804)
  );

  defparam id02327.INIT = 8'h3A;
  LUT3 id02327 (
    .ADR0(id04656),
    .ADR1(id04822),
    .ADR2(id04655),
    .O(id04805)
  );

  defparam id02328.INIT = 4'h6;
  LUT2 id02328 (
    .ADR0(id04801),
    .ADR1(id04802),
    .O(id04806)
  );

  defparam id02329.INIT = 16'h9669;
  LUT4 id02329 (
    .ADR0(id04799),
    .ADR1(id04800),
    .ADR2(id04853),
    .ADR3(id04854),
    .O(id04801)
  );

  defparam id02330.INIT = 8'h35;
  LUT3 id02330 (
    .ADR0(id04820),
    .ADR1(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x0 ),
    .ADR2(id04819),
    .O(id04799)
  );

  defparam id02331.INIT = 4'h9;
  LUT2 id02331 (
    .ADR0(id04851),
    .ADR1(id04852),
    .O(id04800)
  );

  defparam id02332.INIT = 16'h9669;
  LUT4 id02332 (
    .ADR0(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x2 ),
    .O(id04851)
  );

  defparam id02333.INIT = 8'hE8;
  LUT3 id02333 (
    .ADR0(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[23].u_compressor42_cell.x2 ),
    .O(id04852)
  );

  defparam id02334.INIT = 16'h7117;
  LUT4 id02334 (
    .ADR0(id04826),
    .ADR1(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x0 ),
    .ADR2(id04825),
    .ADR3(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x3 ),
    .O(id04853)
  );

  defparam id02335.INIT = 16'h6996;
  LUT4 id02335 (
    .ADR0(id04857),
    .ADR1(id04858),
    .ADR2(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x3 ),
    .O(id04854)
  );

  defparam id02336.INIT = 4'h6;
  LUT2 id02336 (
    .ADR0(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x2 ),
    .O(id04857)
  );

  defparam id02337.INIT = 8'hE8;
  LUT3 id02337 (
    .ADR0(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[29].u_compressor42_cell.x2 ),
    .O(id04858)
  );

  defparam id02338.INIT = 8'hB2;
  LUT3 id02338 (
    .ADR0(id04653),
    .ADR1(id04654),
    .ADR2(id04821),
    .O(id04802)
  );

  defparam id02339.INIT = 8'hB2;
  LUT3 id02339 (
    .ADR0(id04669),
    .ADR1(id04670),
    .ADR2(id04659),
    .O(id04818)
  );

  defparam id02340.INIT = 16'h8E71;
  LUT4 id02340 (
    .ADR0(id04823),
    .ADR1(id04814),
    .ADR2(id04813),
    .ADR3(id04855),
    .O(\net_Buf-pad-result[31] )
  );

  defparam id02341.INIT = 4'h9;
  LUT2 id02341 (
    .ADR0(id04856),
    .ADR1(id04845),
    .O(id04855)
  );

  defparam id02342.INIT = 4'h9;
  LUT2 id02342 (
    .ADR0(id04846),
    .ADR1(id04843),
    .O(id04856)
  );

  defparam id02343.INIT = 8'hC5;
  LUT3 id02343 (
    .ADR0(id04806),
    .ADR1(id04818),
    .ADR2(id04817),
    .O(id04846)
  );

  defparam id02344.INIT = 4'h6;
  LUT2 id02344 (
    .ADR0(id04844),
    .ADR1(id04849),
    .O(id04843)
  );

  defparam id02345.INIT = 16'h9669;
  LUT4 id02345 (
    .ADR0(id04850),
    .ADR1(id04847),
    .ADR2(id04848),
    .ADR3(id04837),
    .O(id04844)
  );

  defparam id02346.INIT = 8'h3A;
  LUT3 id02346 (
    .ADR0(id04804),
    .ADR1(id04808),
    .ADR2(id04803),
    .O(id04850)
  );

  defparam id02347.INIT = 4'h9;
  LUT2 id02347 (
    .ADR0(id04838),
    .ADR1(id04835),
    .O(id04847)
  );

  defparam id02348.INIT = 16'h9669;
  LUT4 id02348 (
    .ADR0(id04836),
    .ADR1(id04841),
    .ADR2(id04842),
    .ADR3(id04839),
    .O(id04838)
  );

  defparam id02349.INIT = 8'h35;
  LUT3 id02349 (
    .ADR0(id04798),
    .ADR1(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x0 ),
    .ADR2(id04797),
    .O(id04836)
  );

  defparam id02350.INIT = 4'h9;
  LUT2 id02350 (
    .ADR0(id04840),
    .ADR1(id04829),
    .O(id04841)
  );

  defparam id02351.INIT = 16'h9669;
  LUT4 id02351 (
    .ADR0(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04840)
  );

  defparam id02352.INIT = 8'hE8;
  LUT3 id02352 (
    .ADR0(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[8].u_compressor42_cell.x2 ),
    .O(id04829)
  );

  defparam id02353.INIT = 16'h7117;
  LUT4 id02353 (
    .ADR0(id04796),
    .ADR1(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x0 ),
    .ADR2(id04795),
    .ADR3(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x3 ),
    .O(id04842)
  );

  defparam id02354.INIT = 16'h6996;
  LUT4 id02354 (
    .ADR0(id04830),
    .ADR1(id04827),
    .ADR2(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x3 ),
    .O(id04839)
  );

  defparam id02355.INIT = 4'h6;
  LUT2 id02355 (
    .ADR0(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04830)
  );

  defparam id02356.INIT = 8'hE8;
  LUT3 id02356 (
    .ADR0(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[16].u_compressor42_cell.x2 ),
    .O(id04827)
  );

  defparam id02357.INIT = 8'h71;
  LUT3 id02357 (
    .ADR0(id04809),
    .ADR1(id04807),
    .ADR2(id04810),
    .O(id04835)
  );

  defparam id02358.INIT = 8'h3A;
  LUT3 id02358 (
    .ADR0(id04802),
    .ADR1(id04854),
    .ADR2(id04801),
    .O(id04848)
  );

  defparam id02359.INIT = 4'h6;
  LUT2 id02359 (
    .ADR0(id04828),
    .ADR1(id04833),
    .O(id04837)
  );

  defparam id02360.INIT = 16'h6996;
  LUT4 id02360 (
    .ADR0(id04834),
    .ADR1(id04831),
    .ADR2(id04832),
    .ADR3(id04771),
    .O(id04828)
  );

  defparam id02361.INIT = 8'h35;
  LUT3 id02361 (
    .ADR0(id04852),
    .ADR1(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x0 ),
    .ADR2(id04851),
    .O(id04834)
  );

  defparam id02362.INIT = 4'h9;
  LUT2 id02362 (
    .ADR0(id04772),
    .ADR1(id04769),
    .O(id04831)
  );

  defparam id02363.INIT = 16'h9669;
  LUT4 id02363 (
    .ADR0(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x2 ),
    .O(id04772)
  );

  defparam id02364.INIT = 8'hE8;
  LUT3 id02364 (
    .ADR0(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_1.CELLS[24].u_compressor42_cell.x2 ),
    .O(id04769)
  );

  defparam id02365.INIT = 16'h7117;
  LUT4 id02365 (
    .ADR0(id04858),
    .ADR1(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x0 ),
    .ADR2(id04857),
    .ADR3(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x3 ),
    .O(id04832)
  );

  defparam id02366.INIT = 16'h6996;
  LUT4 id02366 (
    .ADR0(id04770),
    .ADR1(id04775),
    .ADR2(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x3 ),
    .O(id04771)
  );

  defparam id02367.INIT = 4'h6;
  LUT2 id02367 (
    .ADR0(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[31].u_compressor42_cell.x2 ),
    .O(id04770)
  );

  defparam id02368.INIT = 8'hE8;
  LUT3 id02368 (
    .ADR0(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_0.CELLS[30].u_compressor42_cell.x2 ),
    .O(id04775)
  );

  defparam id02369.INIT = 8'h71;
  LUT3 id02369 (
    .ADR0(id04799),
    .ADR1(id04853),
    .ADR2(id04800),
    .O(id04833)
  );

  defparam id02370.INIT = 8'hB2;
  LUT3 id02370 (
    .ADR0(id04815),
    .ADR1(id04816),
    .ADR2(id04805),
    .O(id04849)
  );

  defparam id02371.INIT = 8'h2B;
  LUT3 id02371 (
    .ADR0(id04811),
    .ADR1(id04812),
    .ADR2(id03943),
    .O(id04845)
  );

  defparam id02372.INIT = 4'h6;
  LUT2 id02372 (
    .ADR0(id04776),
    .ADR1(id04773),
    .O(\net_Buf-pad-result[32] )
  );

  defparam id02373.INIT = 16'h004F;
  LUT4 id02373 (
    .ADR0(id04823),
    .ADR1(id04824),
    .ADR2(id04774),
    .ADR3(id04763),
    .O(id04776)
  );

  defparam id02374.INIT = 4'h4;
  LUT2 id02374 (
    .ADR0(id04856),
    .ADR1(id04845),
    .O(id04763)
  );

  defparam id02375.INIT = 16'hB0BB;
  LUT4 id02375 (
    .ADR0(id04845),
    .ADR1(id04856),
    .ADR2(id04814),
    .ADR3(id04813),
    .O(id04774)
  );

  defparam id02376.INIT = 4'h6;
  LUT2 id02376 (
    .ADR0(id04764),
    .ADR1(id04761),
    .O(id04773)
  );

  defparam id02377.INIT = 4'h4;
  LUT2 id02377 (
    .ADR0(id04846),
    .ADR1(id04843),
    .O(id04764)
  );

  defparam id02378.INIT = 4'h9;
  LUT2 id02378 (
    .ADR0(id04762),
    .ADR1(id04767),
    .O(id04761)
  );

  defparam id02379.INIT = 8'h3A;
  LUT3 id02379 (
    .ADR0(id04849),
    .ADR1(id04837),
    .ADR2(id04844),
    .O(id04762)
  );

  defparam id02380.INIT = 4'h6;
  LUT2 id02380 (
    .ADR0(id04768),
    .ADR1(id04765),
    .O(id04767)
  );

  defparam id02381.INIT = 16'h9669;
  LUT4 id02381 (
    .ADR0(id04766),
    .ADR1(id04755),
    .ADR2(id04756),
    .ADR3(id04753),
    .O(id04768)
  );

  defparam id02382.INIT = 8'h35;
  LUT3 id02382 (
    .ADR0(id04835),
    .ADR1(id04839),
    .ADR2(id04838),
    .O(id04766)
  );

  defparam id02383.INIT = 4'h9;
  LUT2 id02383 (
    .ADR0(id04754),
    .ADR1(id04759),
    .O(id04755)
  );

  defparam id02384.INIT = 16'h6996;
  LUT4 id02384 (
    .ADR0(id04760),
    .ADR1(id04757),
    .ADR2(id04758),
    .ADR3(id04747),
    .O(id04754)
  );

  defparam id02385.INIT = 8'h35;
  LUT3 id02385 (
    .ADR0(id04829),
    .ADR1(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x0 ),
    .ADR2(id04840),
    .O(id04760)
  );

  defparam id02386.INIT = 4'h9;
  LUT2 id02386 (
    .ADR0(id04748),
    .ADR1(id04745),
    .O(id04757)
  );

  defparam id02387.INIT = 16'h9669;
  LUT4 id02387 (
    .ADR0(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_3.CELLS[10].u_compressor42_cell.x2 ),
    .O(id04748)
  );

  defparam id02388.INIT = 8'hE8;
  LUT3 id02388 (
    .ADR0(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_3.CELLS[9].u_compressor42_cell.x2 ),
    .O(id04745)
  );

  defparam id02389.INIT = 16'h7117;
  LUT4 id02389 (
    .ADR0(id04827),
    .ADR1(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x0 ),
    .ADR2(id04830),
    .ADR3(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x3 ),
    .O(id04758)
  );

  defparam id02390.INIT = 16'h6996;
  LUT4 id02390 (
    .ADR0(id04746),
    .ADR1(id04751),
    .ADR2(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x0 ),
    .ADR3(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x3 ),
    .O(id04747)
  );

  defparam id02391.INIT = 4'h6;
  LUT2 id02391 (
    .ADR0(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[18].u_compressor42_cell.x2 ),
    .O(id04746)
  );

  defparam id02392.INIT = 8'hE8;
  LUT3 id02392 (
    .ADR0(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x1 ),
    .ADR1(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x3 ),
    .ADR2(\u_compressor42_l0_2.CELLS[17].u_compressor42_cell.x2 ),
    .O(id04751)
  );

  defparam id02393.INIT = 8'hB2;
  LUT3 id02393 (
    .ADR0(id04836),
    .ADR1(id04841),
    .ADR2(id04842),
    .O(id04759)
  );

  defparam id02394.INIT = 8'h35;
  LUT3 id02394 (
    .ADR0(id04771),
    .ADR1(id04833),
    .ADR2(id04828),
    .O(id04756)
  );

  defparam id02395.INIT = 4'h6;
  LUT2 id02395 (
    .ADR0(id04752),
    .ADR1(id04749),
    .O(id04753)
  );

  defparam id02396.INIT = 16'h9669;
  LUT4 id02396 (
    .ADR0(id04750),
    .ADR1(id04789),
    .ADR2(id04790),
    .ADR3(id04787),
    .O(id04752)
  );

  defparam id02397.INIT = 8'h35;
  LUT3 id02397 (
    .ADR0(id04769),
    .ADR1(\u_compressor42_l0_1.CELLS[25].u_compressor42_cell.x0 ),
    .ADR2(id04772),
    .O(id04750)
  );

  defparam id02398.INIT = 4'h9;
  LUT2 id02398 (
    .ADR0(id04788),
    .ADR1(id04793),
    .O(id04789)
  );

  defparam id02399.INIT = 16'h9669;
  LUT4 id02399 (
    .ADR0(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x0 ),
    .ADR1(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x1 ),
    .ADR2(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x3 ),
    .ADR3(\u_compressor42_l0_1.CELLS[26].u_compressor42_cell.x2 ),
    .O(id04788)
  );

  IBUF \Buf-pad-multiplicand[31]  (
    .I(multiplicand[31]),
    .O(\net_Buf-pad-multiplicand[31] )
  );

  IBUF \Buf-pad-multiplicand[30]  (
    .I(multiplicand[30]),
    .O(\net_Buf-pad-multiplicand[30] )
  );

  IBUF \Buf-pad-multiplicand[29]  (
    .I(multiplicand[29]),
    .O(\net_Buf-pad-multiplicand[29] )
  );

  IBUF \Buf-pad-multiplicand[28]  (
    .I(multiplicand[28]),
    .O(\net_Buf-pad-multiplicand[28] )
  );

  IBUF \Buf-pad-multiplicand[27]  (
    .I(multiplicand[27]),
    .O(\net_Buf-pad-multiplicand[27] )
  );

  IBUF \Buf-pad-multiplicand[26]  (
    .I(multiplicand[26]),
    .O(\net_Buf-pad-multiplicand[26] )
  );

  IBUF \Buf-pad-multiplicand[25]  (
    .I(multiplicand[25]),
    .O(\net_Buf-pad-multiplicand[25] )
  );

  IBUF \Buf-pad-multiplicand[24]  (
    .I(multiplicand[24]),
    .O(\net_Buf-pad-multiplicand[24] )
  );

  IBUF \Buf-pad-multiplicand[23]  (
    .I(multiplicand[23]),
    .O(\net_Buf-pad-multiplicand[23] )
  );

  IBUF \Buf-pad-multiplicand[22]  (
    .I(multiplicand[22]),
    .O(\net_Buf-pad-multiplicand[22] )
  );

  IBUF \Buf-pad-multiplicand[21]  (
    .I(multiplicand[21]),
    .O(\net_Buf-pad-multiplicand[21] )
  );

  IBUF \Buf-pad-multiplicand[20]  (
    .I(multiplicand[20]),
    .O(\net_Buf-pad-multiplicand[20] )
  );

  IBUF \Buf-pad-multiplicand[19]  (
    .I(multiplicand[19]),
    .O(\net_Buf-pad-multiplicand[19] )
  );

  IBUF \Buf-pad-multiplicand[18]  (
    .I(multiplicand[18]),
    .O(\net_Buf-pad-multiplicand[18] )
  );

  IBUF \Buf-pad-multiplicand[17]  (
    .I(multiplicand[17]),
    .O(\net_Buf-pad-multiplicand[17] )
  );

  IBUF \Buf-pad-multiplicand[16]  (
    .I(multiplicand[16]),
    .O(\net_Buf-pad-multiplicand[16] )
  );

  IBUF \Buf-pad-multiplicand[15]  (
    .I(multiplicand[15]),
    .O(\net_Buf-pad-multiplicand[15] )
  );

  IBUF \Buf-pad-multiplicand[14]  (
    .I(multiplicand[14]),
    .O(\net_Buf-pad-multiplicand[14] )
  );

  IBUF \Buf-pad-multiplicand[13]  (
    .I(multiplicand[13]),
    .O(\net_Buf-pad-multiplicand[13] )
  );

  IBUF \Buf-pad-multiplicand[12]  (
    .I(multiplicand[12]),
    .O(\net_Buf-pad-multiplicand[12] )
  );

  IBUF \Buf-pad-multiplicand[11]  (
    .I(multiplicand[11]),
    .O(\net_Buf-pad-multiplicand[11] )
  );

  IBUF \Buf-pad-multiplicand[10]  (
    .I(multiplicand[10]),
    .O(\net_Buf-pad-multiplicand[10] )
  );

  IBUF \Buf-pad-multiplicand[9]  (
    .I(multiplicand[9]),
    .O(\net_Buf-pad-multiplicand[9] )
  );

  IBUF \Buf-pad-multiplicand[8]  (
    .I(multiplicand[8]),
    .O(\net_Buf-pad-multiplicand[8] )
  );

  IBUF \Buf-pad-multiplicand[7]  (
    .I(multiplicand[7]),
    .O(\net_Buf-pad-multiplicand[7] )
  );

  IBUF \Buf-pad-multiplicand[6]  (
    .I(multiplicand[6]),
    .O(\net_Buf-pad-multiplicand[6] )
  );

  IBUF \Buf-pad-multiplicand[5]  (
    .I(multiplicand[5]),
    .O(\net_Buf-pad-multiplicand[5] )
  );

  IBUF \Buf-pad-multiplicand[4]  (
    .I(multiplicand[4]),
    .O(\net_Buf-pad-multiplicand[4] )
  );

  IBUF \Buf-pad-multiplicand[3]  (
    .I(multiplicand[3]),
    .O(\net_Buf-pad-multiplicand[3] )
  );

  IBUF \Buf-pad-multiplicand[2]  (
    .I(multiplicand[2]),
    .O(\net_Buf-pad-multiplicand[2] )
  );

  IBUF \Buf-pad-multiplicand[1]  (
    .I(multiplicand[1]),
    .O(\net_Buf-pad-multiplicand[1] )
  );

  IBUF \Buf-pad-multiplicand[0]  (
    .I(multiplicand[0]),
    .O(\net_Buf-pad-multiplicand[0] )
  );

  IBUF \Buf-pad-multiplier[31]  (
    .I(multiplier[31]),
    .O(\net_Buf-pad-multiplier[31] )
  );

  IBUF \Buf-pad-multiplier[30]  (
    .I(multiplier[30]),
    .O(\net_Buf-pad-multiplier[30] )
  );

  IBUF \Buf-pad-multiplier[29]  (
    .I(multiplier[29]),
    .O(\net_Buf-pad-multiplier[29] )
  );

  IBUF \Buf-pad-multiplier[28]  (
    .I(multiplier[28]),
    .O(\net_Buf-pad-multiplier[28] )
  );

  IBUF \Buf-pad-multiplier[27]  (
    .I(multiplier[27]),
    .O(\net_Buf-pad-multiplier[27] )
  );

  IBUF \Buf-pad-multiplier[26]  (
    .I(multiplier[26]),
    .O(\net_Buf-pad-multiplier[26] )
  );

  IBUF \Buf-pad-multiplier[25]  (
    .I(multiplier[25]),
    .O(\net_Buf-pad-multiplier[25] )
  );

  IBUF \Buf-pad-multiplier[24]  (
    .I(multiplier[24]),
    .O(\net_Buf-pad-multiplier[24] )
  );

  IBUF \Buf-pad-multiplier[23]  (
    .I(multiplier[23]),
    .O(\net_Buf-pad-multiplier[23] )
  );

  IBUF \Buf-pad-multiplier[22]  (
    .I(multiplier[22]),
    .O(\net_Buf-pad-multiplier[22] )
  );

  IBUF \Buf-pad-multiplier[21]  (
    .I(multiplier[21]),
    .O(\net_Buf-pad-multiplier[21] )
  );

  IBUF \Buf-pad-multiplier[20]  (
    .I(multiplier[20]),
    .O(\net_Buf-pad-multiplier[20] )
  );

  IBUF \Buf-pad-multiplier[19]  (
    .I(multiplier[19]),
    .O(\net_Buf-pad-multiplier[19] )
  );

  IBUF \Buf-pad-multiplier[18]  (
    .I(multiplier[18]),
    .O(\net_Buf-pad-multiplier[18] )
  );

  IBUF \Buf-pad-multiplier[17]  (
    .I(multiplier[17]),
    .O(\net_Buf-pad-multiplier[17] )
  );

  IBUF \Buf-pad-multiplier[16]  (
    .I(multiplier[16]),
    .O(\net_Buf-pad-multiplier[16] )
  );

  IBUF \Buf-pad-multiplier[15]  (
    .I(multiplier[15]),
    .O(\net_Buf-pad-multiplier[15] )
  );

  IBUF \Buf-pad-multiplier[14]  (
    .I(multiplier[14]),
    .O(\net_Buf-pad-multiplier[14] )
  );

  IBUF \Buf-pad-multiplier[13]  (
    .I(multiplier[13]),
    .O(\net_Buf-pad-multiplier[13] )
  );

  IBUF \Buf-pad-multiplier[12]  (
    .I(multiplier[12]),
    .O(\net_Buf-pad-multiplier[12] )
  );

  IBUF \Buf-pad-multiplier[11]  (
    .I(multiplier[11]),
    .O(\net_Buf-pad-multiplier[11] )
  );

  IBUF \Buf-pad-multiplier[10]  (
    .I(multiplier[10]),
    .O(\net_Buf-pad-multiplier[10] )
  );

  IBUF \Buf-pad-multiplier[9]  (
    .I(multiplier[9]),
    .O(\net_Buf-pad-multiplier[9] )
  );

  IBUF \Buf-pad-multiplier[8]  (
    .I(multiplier[8]),
    .O(\net_Buf-pad-multiplier[8] )
  );

  IBUF \Buf-pad-multiplier[7]  (
    .I(multiplier[7]),
    .O(\net_Buf-pad-multiplier[7] )
  );

  IBUF \Buf-pad-multiplier[6]  (
    .I(multiplier[6]),
    .O(\net_Buf-pad-multiplier[6] )
  );

  IBUF \Buf-pad-multiplier[5]  (
    .I(multiplier[5]),
    .O(\net_Buf-pad-multiplier[5] )
  );

  IBUF \Buf-pad-multiplier[4]  (
    .I(multiplier[4]),
    .O(\net_Buf-pad-multiplier[4] )
  );

  IBUF \Buf-pad-multiplier[3]  (
    .I(multiplier[3]),
    .O(\net_Buf-pad-multiplier[3] )
  );

  IBUF \Buf-pad-multiplier[2]  (
    .I(multiplier[2]),
    .O(\net_Buf-pad-multiplier[2] )
  );

  IBUF \Buf-pad-multiplier[1]  (
    .I(multiplier[1]),
    .O(\net_Buf-pad-multiplier[1] )
  );

  IBUF \Buf-pad-multiplier[0]  (
    .I(multiplier[0]),
    .O(\net_Buf-pad-multiplier[0] )
  );

  IPAD \multiplicand[31]_ipad  (
    .PAD(multiplicand[31])
  );

  IPAD \multiplicand[30]_ipad  (
    .PAD(multiplicand[30])
  );

  IPAD \multiplicand[29]_ipad  (
    .PAD(multiplicand[29])
  );

  IPAD \multiplicand[28]_ipad  (
    .PAD(multiplicand[28])
  );

  IPAD \multiplicand[27]_ipad  (
    .PAD(multiplicand[27])
  );

  IPAD \multiplicand[26]_ipad  (
    .PAD(multiplicand[26])
  );

  IPAD \multiplicand[25]_ipad  (
    .PAD(multiplicand[25])
  );

  IPAD \multiplicand[24]_ipad  (
    .PAD(multiplicand[24])
  );

  IPAD \multiplicand[23]_ipad  (
    .PAD(multiplicand[23])
  );

  IPAD \multiplicand[22]_ipad  (
    .PAD(multiplicand[22])
  );

  IPAD \multiplicand[21]_ipad  (
    .PAD(multiplicand[21])
  );

  IPAD \multiplicand[20]_ipad  (
    .PAD(multiplicand[20])
  );

  IPAD \multiplicand[19]_ipad  (
    .PAD(multiplicand[19])
  );

  IPAD \multiplicand[18]_ipad  (
    .PAD(multiplicand[18])
  );

  IPAD \multiplicand[17]_ipad  (
    .PAD(multiplicand[17])
  );

  IPAD \multiplicand[16]_ipad  (
    .PAD(multiplicand[16])
  );

  IPAD \multiplicand[15]_ipad  (
    .PAD(multiplicand[15])
  );

  IPAD \multiplicand[14]_ipad  (
    .PAD(multiplicand[14])
  );

  IPAD \multiplicand[13]_ipad  (
    .PAD(multiplicand[13])
  );

  IPAD \multiplicand[12]_ipad  (
    .PAD(multiplicand[12])
  );

  IPAD \multiplicand[11]_ipad  (
    .PAD(multiplicand[11])
  );

  IPAD \multiplicand[10]_ipad  (
    .PAD(multiplicand[10])
  );

  IPAD \multiplicand[9]_ipad  (
    .PAD(multiplicand[9])
  );

  IPAD \multiplicand[8]_ipad  (
    .PAD(multiplicand[8])
  );

  IPAD \multiplicand[7]_ipad  (
    .PAD(multiplicand[7])
  );

  IPAD \multiplicand[6]_ipad  (
    .PAD(multiplicand[6])
  );

  IPAD \multiplicand[5]_ipad  (
    .PAD(multiplicand[5])
  );

  IPAD \multiplicand[4]_ipad  (
    .PAD(multiplicand[4])
  );

  IPAD \multiplicand[3]_ipad  (
    .PAD(multiplicand[3])
  );

  IPAD \multiplicand[2]_ipad  (
    .PAD(multiplicand[2])
  );

  IPAD \multiplicand[1]_ipad  (
    .PAD(multiplicand[1])
  );

  IPAD \multiplicand[0]_ipad  (
    .PAD(multiplicand[0])
  );

  IPAD \multiplier[31]_ipad  (
    .PAD(multiplier[31])
  );

  IPAD \multiplier[30]_ipad  (
    .PAD(multiplier[30])
  );

  IPAD \multiplier[29]_ipad  (
    .PAD(multiplier[29])
  );

  IPAD \multiplier[28]_ipad  (
    .PAD(multiplier[28])
  );

  IPAD \multiplier[27]_ipad  (
    .PAD(multiplier[27])
  );

  IPAD \multiplier[26]_ipad  (
    .PAD(multiplier[26])
  );

  IPAD \multiplier[25]_ipad  (
    .PAD(multiplier[25])
  );

  IPAD \multiplier[24]_ipad  (
    .PAD(multiplier[24])
  );

  IPAD \multiplier[23]_ipad  (
    .PAD(multiplier[23])
  );

  IPAD \multiplier[22]_ipad  (
    .PAD(multiplier[22])
  );

  IPAD \multiplier[21]_ipad  (
    .PAD(multiplier[21])
  );

  IPAD \multiplier[20]_ipad  (
    .PAD(multiplier[20])
  );

  IPAD \multiplier[19]_ipad  (
    .PAD(multiplier[19])
  );

  IPAD \multiplier[18]_ipad  (
    .PAD(multiplier[18])
  );

  IPAD \multiplier[17]_ipad  (
    .PAD(multiplier[17])
  );

  IPAD \multiplier[16]_ipad  (
    .PAD(multiplier[16])
  );

  IPAD \multiplier[15]_ipad  (
    .PAD(multiplier[15])
  );

  IPAD \multiplier[14]_ipad  (
    .PAD(multiplier[14])
  );

  IPAD \multiplier[13]_ipad  (
    .PAD(multiplier[13])
  );

  IPAD \multiplier[12]_ipad  (
    .PAD(multiplier[12])
  );

  IPAD \multiplier[11]_ipad  (
    .PAD(multiplier[11])
  );

  IPAD \multiplier[10]_ipad  (
    .PAD(multiplier[10])
  );

  IPAD \multiplier[9]_ipad  (
    .PAD(multiplier[9])
  );

  IPAD \multiplier[8]_ipad  (
    .PAD(multiplier[8])
  );

  IPAD \multiplier[7]_ipad  (
    .PAD(multiplier[7])
  );

  IPAD \multiplier[6]_ipad  (
    .PAD(multiplier[6])
  );

  IPAD \multiplier[5]_ipad  (
    .PAD(multiplier[5])
  );

  IPAD \multiplier[4]_ipad  (
    .PAD(multiplier[4])
  );

  IPAD \multiplier[3]_ipad  (
    .PAD(multiplier[3])
  );

  IPAD \multiplier[2]_ipad  (
    .PAD(multiplier[2])
  );

  IPAD \multiplier[1]_ipad  (
    .PAD(multiplier[1])
  );

  IPAD \multiplier[0]_ipad  (
    .PAD(multiplier[0])
  );

  OBUF \Buf-pad-result[63]  (
    .I(\net_Buf-pad-result[63] ),
    .O(result[63])
  );

  OBUF \Buf-pad-result[62]  (
    .I(\net_Buf-pad-result[62] ),
    .O(result[62])
  );

  OBUF \Buf-pad-result[61]  (
    .I(\net_Buf-pad-result[61] ),
    .O(result[61])
  );

  OBUF \Buf-pad-result[60]  (
    .I(\net_Buf-pad-result[60] ),
    .O(result[60])
  );

  OBUF \Buf-pad-result[59]  (
    .I(\net_Buf-pad-result[59] ),
    .O(result[59])
  );

  OBUF \Buf-pad-result[58]  (
    .I(\net_Buf-pad-result[58] ),
    .O(result[58])
  );

  OBUF \Buf-pad-result[57]  (
    .I(\net_Buf-pad-result[57] ),
    .O(result[57])
  );

  OBUF \Buf-pad-result[56]  (
    .I(\net_Buf-pad-result[56] ),
    .O(result[56])
  );

  OBUF \Buf-pad-result[55]  (
    .I(\net_Buf-pad-result[55] ),
    .O(result[55])
  );

  OBUF \Buf-pad-result[54]  (
    .I(\net_Buf-pad-result[54] ),
    .O(result[54])
  );

  OBUF \Buf-pad-result[53]  (
    .I(\net_Buf-pad-result[53] ),
    .O(result[53])
  );

  OBUF \Buf-pad-result[52]  (
    .I(\net_Buf-pad-result[52] ),
    .O(result[52])
  );

  OBUF \Buf-pad-result[51]  (
    .I(\net_Buf-pad-result[51] ),
    .O(result[51])
  );

  OBUF \Buf-pad-result[50]  (
    .I(\net_Buf-pad-result[50] ),
    .O(result[50])
  );

  OBUF \Buf-pad-result[49]  (
    .I(\net_Buf-pad-result[49] ),
    .O(result[49])
  );

  OBUF \Buf-pad-result[48]  (
    .I(\net_Buf-pad-result[48] ),
    .O(result[48])
  );

  OBUF \Buf-pad-result[47]  (
    .I(\net_Buf-pad-result[47] ),
    .O(result[47])
  );

  OBUF \Buf-pad-result[46]  (
    .I(\net_Buf-pad-result[46] ),
    .O(result[46])
  );

  OBUF \Buf-pad-result[45]  (
    .I(\net_Buf-pad-result[45] ),
    .O(result[45])
  );

  OBUF \Buf-pad-result[44]  (
    .I(\net_Buf-pad-result[44] ),
    .O(result[44])
  );

  OBUF \Buf-pad-result[43]  (
    .I(\net_Buf-pad-result[43] ),
    .O(result[43])
  );

  OBUF \Buf-pad-result[42]  (
    .I(\net_Buf-pad-result[42] ),
    .O(result[42])
  );

  OBUF \Buf-pad-result[41]  (
    .I(\net_Buf-pad-result[41] ),
    .O(result[41])
  );

  OBUF \Buf-pad-result[40]  (
    .I(\net_Buf-pad-result[40] ),
    .O(result[40])
  );

  OBUF \Buf-pad-result[39]  (
    .I(\net_Buf-pad-result[39] ),
    .O(result[39])
  );

  OBUF \Buf-pad-result[38]  (
    .I(\net_Buf-pad-result[38] ),
    .O(result[38])
  );

  OBUF \Buf-pad-result[37]  (
    .I(\net_Buf-pad-result[37] ),
    .O(result[37])
  );

  OBUF \Buf-pad-result[36]  (
    .I(\net_Buf-pad-result[36] ),
    .O(result[36])
  );

  OBUF \Buf-pad-result[35]  (
    .I(\net_Buf-pad-result[35] ),
    .O(result[35])
  );

  OBUF \Buf-pad-result[34]  (
    .I(\net_Buf-pad-result[34] ),
    .O(result[34])
  );

  OBUF \Buf-pad-result[33]  (
    .I(\net_Buf-pad-result[33] ),
    .O(result[33])
  );

  OBUF \Buf-pad-result[32]  (
    .I(\net_Buf-pad-result[32] ),
    .O(result[32])
  );

  OBUF \Buf-pad-result[31]  (
    .I(\net_Buf-pad-result[31] ),
    .O(result[31])
  );

  OBUF \Buf-pad-result[30]  (
    .I(\net_Buf-pad-result[30] ),
    .O(result[30])
  );

  OBUF \Buf-pad-result[29]  (
    .I(\net_Buf-pad-result[29] ),
    .O(result[29])
  );

  OBUF \Buf-pad-result[28]  (
    .I(\net_Buf-pad-result[28] ),
    .O(result[28])
  );

  OBUF \Buf-pad-result[27]  (
    .I(\net_Buf-pad-result[27] ),
    .O(result[27])
  );

  OBUF \Buf-pad-result[26]  (
    .I(\net_Buf-pad-result[26] ),
    .O(result[26])
  );

  OBUF \Buf-pad-result[25]  (
    .I(\net_Buf-pad-result[25] ),
    .O(result[25])
  );

  OBUF \Buf-pad-result[24]  (
    .I(\net_Buf-pad-result[24] ),
    .O(result[24])
  );

  OBUF \Buf-pad-result[23]  (
    .I(\net_Buf-pad-result[23] ),
    .O(result[23])
  );

  OBUF \Buf-pad-result[22]  (
    .I(\net_Buf-pad-result[22] ),
    .O(result[22])
  );

  OBUF \Buf-pad-result[21]  (
    .I(\net_Buf-pad-result[21] ),
    .O(result[21])
  );

  OBUF \Buf-pad-result[20]  (
    .I(\net_Buf-pad-result[20] ),
    .O(result[20])
  );

  OBUF \Buf-pad-result[19]  (
    .I(\net_Buf-pad-result[19] ),
    .O(result[19])
  );

  OBUF \Buf-pad-result[18]  (
    .I(\net_Buf-pad-result[18] ),
    .O(result[18])
  );

  OBUF \Buf-pad-result[17]  (
    .I(\net_Buf-pad-result[17] ),
    .O(result[17])
  );

  OBUF \Buf-pad-result[16]  (
    .I(\net_Buf-pad-result[16] ),
    .O(result[16])
  );

  OBUF \Buf-pad-result[15]  (
    .I(\net_Buf-pad-result[15] ),
    .O(result[15])
  );

  OBUF \Buf-pad-result[14]  (
    .I(\net_Buf-pad-result[14] ),
    .O(result[14])
  );

  OBUF \Buf-pad-result[13]  (
    .I(\net_Buf-pad-result[13] ),
    .O(result[13])
  );

  OBUF \Buf-pad-result[12]  (
    .I(\net_Buf-pad-result[12] ),
    .O(result[12])
  );

  OBUF \Buf-pad-result[11]  (
    .I(\net_Buf-pad-result[11] ),
    .O(result[11])
  );

  OBUF \Buf-pad-result[10]  (
    .I(\net_Buf-pad-result[10] ),
    .O(result[10])
  );

  OBUF \Buf-pad-result[9]  (
    .I(\net_Buf-pad-result[9] ),
    .O(result[9])
  );

  OBUF \Buf-pad-result[8]  (
    .I(\net_Buf-pad-result[8] ),
    .O(result[8])
  );

  OBUF \Buf-pad-result[7]  (
    .I(\net_Buf-pad-result[7] ),
    .O(result[7])
  );

  OBUF \Buf-pad-result[6]  (
    .I(\net_Buf-pad-result[6] ),
    .O(result[6])
  );

  OBUF \Buf-pad-result[5]  (
    .I(\net_Buf-pad-result[5] ),
    .O(result[5])
  );

  OBUF \Buf-pad-result[4]  (
    .I(\net_Buf-pad-result[4] ),
    .O(result[4])
  );

  OBUF \Buf-pad-result[3]  (
    .I(\net_Buf-pad-result[3] ),
    .O(result[3])
  );

  OBUF \Buf-pad-result[2]  (
    .I(\net_Buf-pad-result[2] ),
    .O(result[2])
  );

  OBUF \Buf-pad-result[1]  (
    .I(\net_Buf-pad-result[1] ),
    .O(result[1])
  );

  OBUF \Buf-pad-result[0]  (
    .I(\net_Buf-pad-result[0] ),
    .O(result[0])
  );

  OPAD \result[63]_opad  (
    .PAD(result[63])
  );

  OPAD \result[62]_opad  (
    .PAD(result[62])
  );

  OPAD \result[61]_opad  (
    .PAD(result[61])
  );

  OPAD \result[60]_opad  (
    .PAD(result[60])
  );

  OPAD \result[59]_opad  (
    .PAD(result[59])
  );

  OPAD \result[58]_opad  (
    .PAD(result[58])
  );

  OPAD \result[57]_opad  (
    .PAD(result[57])
  );

  OPAD \result[56]_opad  (
    .PAD(result[56])
  );

  OPAD \result[55]_opad  (
    .PAD(result[55])
  );

  OPAD \result[54]_opad  (
    .PAD(result[54])
  );

  OPAD \result[53]_opad  (
    .PAD(result[53])
  );

  OPAD \result[52]_opad  (
    .PAD(result[52])
  );

  OPAD \result[51]_opad  (
    .PAD(result[51])
  );

  OPAD \result[50]_opad  (
    .PAD(result[50])
  );

  OPAD \result[49]_opad  (
    .PAD(result[49])
  );

  OPAD \result[48]_opad  (
    .PAD(result[48])
  );

  OPAD \result[47]_opad  (
    .PAD(result[47])
  );

  OPAD \result[46]_opad  (
    .PAD(result[46])
  );

  OPAD \result[45]_opad  (
    .PAD(result[45])
  );

  OPAD \result[44]_opad  (
    .PAD(result[44])
  );

  OPAD \result[43]_opad  (
    .PAD(result[43])
  );

  OPAD \result[42]_opad  (
    .PAD(result[42])
  );

  OPAD \result[41]_opad  (
    .PAD(result[41])
  );

  OPAD \result[40]_opad  (
    .PAD(result[40])
  );

  OPAD \result[39]_opad  (
    .PAD(result[39])
  );

  OPAD \result[38]_opad  (
    .PAD(result[38])
  );

  OPAD \result[37]_opad  (
    .PAD(result[37])
  );

  OPAD \result[36]_opad  (
    .PAD(result[36])
  );

  OPAD \result[35]_opad  (
    .PAD(result[35])
  );

  OPAD \result[34]_opad  (
    .PAD(result[34])
  );

  OPAD \result[33]_opad  (
    .PAD(result[33])
  );

  OPAD \result[32]_opad  (
    .PAD(result[32])
  );

  OPAD \result[31]_opad  (
    .PAD(result[31])
  );

  OPAD \result[30]_opad  (
    .PAD(result[30])
  );

  OPAD \result[29]_opad  (
    .PAD(result[29])
  );

  OPAD \result[28]_opad  (
    .PAD(result[28])
  );

  OPAD \result[27]_opad  (
    .PAD(result[27])
  );

  OPAD \result[26]_opad  (
    .PAD(result[26])
  );

  OPAD \result[25]_opad  (
    .PAD(result[25])
  );

  OPAD \result[24]_opad  (
    .PAD(result[24])
  );

  OPAD \result[23]_opad  (
    .PAD(result[23])
  );

  OPAD \result[22]_opad  (
    .PAD(result[22])
  );

  OPAD \result[21]_opad  (
    .PAD(result[21])
  );

  OPAD \result[20]_opad  (
    .PAD(result[20])
  );

  OPAD \result[19]_opad  (
    .PAD(result[19])
  );

  OPAD \result[18]_opad  (
    .PAD(result[18])
  );

  OPAD \result[17]_opad  (
    .PAD(result[17])
  );

  OPAD \result[16]_opad  (
    .PAD(result[16])
  );

  OPAD \result[15]_opad  (
    .PAD(result[15])
  );

  OPAD \result[14]_opad  (
    .PAD(result[14])
  );

  OPAD \result[13]_opad  (
    .PAD(result[13])
  );

  OPAD \result[12]_opad  (
    .PAD(result[12])
  );

  OPAD \result[11]_opad  (
    .PAD(result[11])
  );

  OPAD \result[10]_opad  (
    .PAD(result[10])
  );

  OPAD \result[9]_opad  (
    .PAD(result[9])
  );

  OPAD \result[8]_opad  (
    .PAD(result[8])
  );

  OPAD \result[7]_opad  (
    .PAD(result[7])
  );

  OPAD \result[6]_opad  (
    .PAD(result[6])
  );

  OPAD \result[5]_opad  (
    .PAD(result[5])
  );

  OPAD \result[4]_opad  (
    .PAD(result[4])
  );

  OPAD \result[3]_opad  (
    .PAD(result[3])
  );

  OPAD \result[2]_opad  (
    .PAD(result[2])
  );

  OPAD \result[1]_opad  (
    .PAD(result[1])
  );

  OPAD \result[0]_opad  (
    .PAD(result[0])
  );

  LOGIC_1 VCC (
    .LOGIC_1_PIN(VCC_NET)
  );

  LOGIC_0 GND (
    .LOGIC_0_PIN(GND_NET)
  );
endmodule
